
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);




    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_keygen.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_keygen.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_keygen.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.grp_process_block_111_112_fu_512.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.grp_process_block_111_112_fu_512.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.grp_process_block_111_112_fu_512.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_keygen.grp_fpr_of_fu_1317.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_keygen.grp_fpr_of_fu_1317.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_keygen.grp_fpr_of_fu_1317.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_keygen.grp_FFT_fu_1324.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_keygen.grp_FFT_fu_1324.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_keygen.grp_FFT_fu_1324.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;
    nodf_module_intf module_intf_7(clock,reset);
    assign module_intf_7.ap_start = AESL_inst_keygen.grp_FFT_fu_1331.ap_start;
    assign module_intf_7.ap_ready = AESL_inst_keygen.grp_FFT_fu_1331.ap_ready;
    assign module_intf_7.ap_done = AESL_inst_keygen.grp_FFT_fu_1331.ap_done;
    assign module_intf_7.ap_continue = 1'b1;
    assign module_intf_7.finish = finish;
    csv_file_dump mstatus_csv_dumper_7;
    nodf_module_monitor module_monitor_7;
    nodf_module_intf module_intf_8(clock,reset);
    assign module_intf_8.ap_start = AESL_inst_keygen.grp_iFFT_fu_1338.ap_start;
    assign module_intf_8.ap_ready = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ready;
    assign module_intf_8.ap_done = AESL_inst_keygen.grp_iFFT_fu_1338.ap_done;
    assign module_intf_8.ap_continue = 1'b1;
    assign module_intf_8.finish = finish;
    csv_file_dump mstatus_csv_dumper_8;
    nodf_module_monitor module_monitor_8;
    nodf_module_intf module_intf_9(clock,reset);
    assign module_intf_9.ap_start = AESL_inst_keygen.grp_iFFT_fu_1345.ap_start;
    assign module_intf_9.ap_ready = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ready;
    assign module_intf_9.ap_done = AESL_inst_keygen.grp_iFFT_fu_1345.ap_done;
    assign module_intf_9.ap_continue = 1'b1;
    assign module_intf_9.finish = finish;
    csv_file_dump mstatus_csv_dumper_9;
    nodf_module_monitor module_monitor_9;
    nodf_module_intf module_intf_10(clock,reset);
    assign module_intf_10.ap_start = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_start;
    assign module_intf_10.ap_ready = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ready;
    assign module_intf_10.ap_done = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_done;
    assign module_intf_10.ap_continue = 1'b1;
    assign module_intf_10.finish = finish;
    csv_file_dump mstatus_csv_dumper_10;
    nodf_module_monitor module_monitor_10;
    nodf_module_intf module_intf_11(clock,reset);
    assign module_intf_11.ap_start = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_start;
    assign module_intf_11.ap_ready = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ready;
    assign module_intf_11.ap_done = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_done;
    assign module_intf_11.ap_continue = 1'b1;
    assign module_intf_11.finish = finish;
    csv_file_dump mstatus_csv_dumper_11;
    nodf_module_monitor module_monitor_11;
    nodf_module_intf module_intf_12(clock,reset);
    assign module_intf_12.ap_start = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_start;
    assign module_intf_12.ap_ready = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ready;
    assign module_intf_12.ap_done = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_done;
    assign module_intf_12.ap_continue = 1'b1;
    assign module_intf_12.finish = finish;
    csv_file_dump mstatus_csv_dumper_12;
    nodf_module_monitor module_monitor_12;
    nodf_module_intf module_intf_13(clock,reset);
    assign module_intf_13.ap_start = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_montysqr_fu_336.ap_start;
    assign module_intf_13.ap_ready = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_montysqr_fu_336.ap_ready;
    assign module_intf_13.ap_done = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_montysqr_fu_336.ap_done;
    assign module_intf_13.ap_continue = 1'b1;
    assign module_intf_13.finish = finish;
    csv_file_dump mstatus_csv_dumper_13;
    nodf_module_monitor module_monitor_13;
    nodf_module_intf module_intf_14(clock,reset);
    assign module_intf_14.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_start;
    assign module_intf_14.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ready;
    assign module_intf_14.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_done;
    assign module_intf_14.ap_continue = 1'b1;
    assign module_intf_14.finish = finish;
    csv_file_dump mstatus_csv_dumper_14;
    nodf_module_monitor module_monitor_14;
    nodf_module_intf module_intf_15(clock,reset);
    assign module_intf_15.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_start;
    assign module_intf_15.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ready;
    assign module_intf_15.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_done;
    assign module_intf_15.ap_continue = 1'b1;
    assign module_intf_15.finish = finish;
    csv_file_dump mstatus_csv_dumper_15;
    nodf_module_monitor module_monitor_15;
    nodf_module_intf module_intf_16(clock,reset);
    assign module_intf_16.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_start;
    assign module_intf_16.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ready;
    assign module_intf_16.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_done;
    assign module_intf_16.ap_continue = 1'b1;
    assign module_intf_16.finish = finish;
    csv_file_dump mstatus_csv_dumper_16;
    nodf_module_monitor module_monitor_16;
    nodf_module_intf module_intf_17(clock,reset);
    assign module_intf_17.ap_start = 1'b0;
    assign module_intf_17.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.grp_modp_montymul_fu_184.ap_ready;
    assign module_intf_17.ap_done = 1'b0;
    assign module_intf_17.ap_continue = 1'b0;
    assign module_intf_17.finish = finish;
    csv_file_dump mstatus_csv_dumper_17;
    nodf_module_monitor module_monitor_17;
    nodf_module_intf module_intf_18(clock,reset);
    assign module_intf_18.ap_start = 1'b0;
    assign module_intf_18.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.grp_modp_montymul_fu_192.ap_ready;
    assign module_intf_18.ap_done = 1'b0;
    assign module_intf_18.ap_continue = 1'b0;
    assign module_intf_18.finish = finish;
    csv_file_dump mstatus_csv_dumper_18;
    nodf_module_monitor module_monitor_18;
    nodf_module_intf module_intf_19(clock,reset);
    assign module_intf_19.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_start;
    assign module_intf_19.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ready;
    assign module_intf_19.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_done;
    assign module_intf_19.ap_continue = 1'b1;
    assign module_intf_19.finish = finish;
    csv_file_dump mstatus_csv_dumper_19;
    nodf_module_monitor module_monitor_19;
    nodf_module_intf module_intf_20(clock,reset);
    assign module_intf_20.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_start;
    assign module_intf_20.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ready;
    assign module_intf_20.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_done;
    assign module_intf_20.ap_continue = 1'b1;
    assign module_intf_20.finish = finish;
    csv_file_dump mstatus_csv_dumper_20;
    nodf_module_monitor module_monitor_20;
    nodf_module_intf module_intf_21(clock,reset);
    assign module_intf_21.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_start;
    assign module_intf_21.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ready;
    assign module_intf_21.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_done;
    assign module_intf_21.ap_continue = 1'b1;
    assign module_intf_21.finish = finish;
    csv_file_dump mstatus_csv_dumper_21;
    nodf_module_monitor module_monitor_21;
    nodf_module_intf module_intf_22(clock,reset);
    assign module_intf_22.ap_start = 1'b0;
    assign module_intf_22.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.grp_modp_montymul_fu_442.ap_ready;
    assign module_intf_22.ap_done = 1'b0;
    assign module_intf_22.ap_continue = 1'b0;
    assign module_intf_22.finish = finish;
    csv_file_dump mstatus_csv_dumper_22;
    nodf_module_monitor module_monitor_22;
    nodf_module_intf module_intf_23(clock,reset);
    assign module_intf_23.ap_start = 1'b0;
    assign module_intf_23.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.grp_modp_montymul_fu_450.ap_ready;
    assign module_intf_23.ap_done = 1'b0;
    assign module_intf_23.ap_continue = 1'b0;
    assign module_intf_23.finish = finish;
    csv_file_dump mstatus_csv_dumper_23;
    nodf_module_monitor module_monitor_23;
    nodf_module_intf module_intf_24(clock,reset);
    assign module_intf_24.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_start;
    assign module_intf_24.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ready;
    assign module_intf_24.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_done;
    assign module_intf_24.ap_continue = 1'b1;
    assign module_intf_24.finish = finish;
    csv_file_dump mstatus_csv_dumper_24;
    nodf_module_monitor module_monitor_24;
    nodf_module_intf module_intf_25(clock,reset);
    assign module_intf_25.ap_start = 1'b0;
    assign module_intf_25.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.grp_modp_montymul_fu_184.ap_ready;
    assign module_intf_25.ap_done = 1'b0;
    assign module_intf_25.ap_continue = 1'b0;
    assign module_intf_25.finish = finish;
    csv_file_dump mstatus_csv_dumper_25;
    nodf_module_monitor module_monitor_25;
    nodf_module_intf module_intf_26(clock,reset);
    assign module_intf_26.ap_start = 1'b0;
    assign module_intf_26.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.grp_modp_montymul_fu_192.ap_ready;
    assign module_intf_26.ap_done = 1'b0;
    assign module_intf_26.ap_continue = 1'b0;
    assign module_intf_26.finish = finish;
    csv_file_dump mstatus_csv_dumper_26;
    nodf_module_monitor module_monitor_26;
    nodf_module_intf module_intf_27(clock,reset);
    assign module_intf_27.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_start;
    assign module_intf_27.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ready;
    assign module_intf_27.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_done;
    assign module_intf_27.ap_continue = 1'b1;
    assign module_intf_27.finish = finish;
    csv_file_dump mstatus_csv_dumper_27;
    nodf_module_monitor module_monitor_27;
    nodf_module_intf module_intf_28(clock,reset);
    assign module_intf_28.ap_start = 1'b0;
    assign module_intf_28.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.y_modp_montymul_fu_200.ap_ready;
    assign module_intf_28.ap_done = 1'b0;
    assign module_intf_28.ap_continue = 1'b0;
    assign module_intf_28.finish = finish;
    csv_file_dump mstatus_csv_dumper_28;
    nodf_module_monitor module_monitor_28;
    nodf_module_intf module_intf_29(clock,reset);
    assign module_intf_29.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_start;
    assign module_intf_29.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ready;
    assign module_intf_29.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_done;
    assign module_intf_29.ap_continue = 1'b1;
    assign module_intf_29.finish = finish;
    csv_file_dump mstatus_csv_dumper_29;
    nodf_module_monitor module_monitor_29;
    nodf_module_intf module_intf_30(clock,reset);
    assign module_intf_30.ap_start = 1'b0;
    assign module_intf_30.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_montymul_fu_255.ap_ready;
    assign module_intf_30.ap_done = 1'b0;
    assign module_intf_30.ap_continue = 1'b0;
    assign module_intf_30.finish = finish;
    csv_file_dump mstatus_csv_dumper_30;
    nodf_module_monitor module_monitor_30;
    nodf_module_intf module_intf_31(clock,reset);
    assign module_intf_31.ap_start = 1'b0;
    assign module_intf_31.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_montymul_fu_265.ap_ready;
    assign module_intf_31.ap_done = 1'b0;
    assign module_intf_31.ap_continue = 1'b0;
    assign module_intf_31.finish = finish;
    csv_file_dump mstatus_csv_dumper_31;
    nodf_module_monitor module_monitor_31;
    nodf_module_intf module_intf_32(clock,reset);
    assign module_intf_32.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_start;
    assign module_intf_32.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ready;
    assign module_intf_32.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_done;
    assign module_intf_32.ap_continue = 1'b1;
    assign module_intf_32.finish = finish;
    csv_file_dump mstatus_csv_dumper_32;
    nodf_module_monitor module_monitor_32;
    nodf_module_intf module_intf_33(clock,reset);
    assign module_intf_33.ap_start = 1'b0;
    assign module_intf_33.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.y_modp_montymul_fu_200.ap_ready;
    assign module_intf_33.ap_done = 1'b0;
    assign module_intf_33.ap_continue = 1'b0;
    assign module_intf_33.finish = finish;
    csv_file_dump mstatus_csv_dumper_33;
    nodf_module_monitor module_monitor_33;
    nodf_module_intf module_intf_34(clock,reset);
    assign module_intf_34.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_start;
    assign module_intf_34.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ready;
    assign module_intf_34.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_done;
    assign module_intf_34.ap_continue = 1'b1;
    assign module_intf_34.finish = finish;
    csv_file_dump mstatus_csv_dumper_34;
    nodf_module_monitor module_monitor_34;
    nodf_module_intf module_intf_35(clock,reset);
    assign module_intf_35.ap_start = 1'b0;
    assign module_intf_35.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.y_modp_montymul_fu_200.ap_ready;
    assign module_intf_35.ap_done = 1'b0;
    assign module_intf_35.ap_continue = 1'b0;
    assign module_intf_35.finish = finish;
    csv_file_dump mstatus_csv_dumper_35;
    nodf_module_monitor module_monitor_35;
    nodf_module_intf module_intf_36(clock,reset);
    assign module_intf_36.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_start;
    assign module_intf_36.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ready;
    assign module_intf_36.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_done;
    assign module_intf_36.ap_continue = 1'b1;
    assign module_intf_36.finish = finish;
    csv_file_dump mstatus_csv_dumper_36;
    nodf_module_monitor module_monitor_36;
    nodf_module_intf module_intf_37(clock,reset);
    assign module_intf_37.ap_start = 1'b0;
    assign module_intf_37.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_montymul_fu_3413.ap_ready;
    assign module_intf_37.ap_done = 1'b0;
    assign module_intf_37.ap_continue = 1'b0;
    assign module_intf_37.finish = finish;
    csv_file_dump mstatus_csv_dumper_37;
    nodf_module_monitor module_monitor_37;
    nodf_module_intf module_intf_38(clock,reset);
    assign module_intf_38.ap_start = 1'b0;
    assign module_intf_38.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_montymul_fu_3425.ap_ready;
    assign module_intf_38.ap_done = 1'b0;
    assign module_intf_38.ap_continue = 1'b0;
    assign module_intf_38.finish = finish;
    csv_file_dump mstatus_csv_dumper_38;
    nodf_module_monitor module_monitor_38;
    nodf_module_intf module_intf_39(clock,reset);
    assign module_intf_39.ap_start = 1'b0;
    assign module_intf_39.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_montymul_fu_3437.ap_ready;
    assign module_intf_39.ap_done = 1'b0;
    assign module_intf_39.ap_continue = 1'b0;
    assign module_intf_39.finish = finish;
    csv_file_dump mstatus_csv_dumper_39;
    nodf_module_monitor module_monitor_39;
    nodf_module_intf module_intf_40(clock,reset);
    assign module_intf_40.ap_start = 1'b0;
    assign module_intf_40.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_montymul_fu_3463.ap_ready;
    assign module_intf_40.ap_done = 1'b0;
    assign module_intf_40.ap_continue = 1'b0;
    assign module_intf_40.finish = finish;
    csv_file_dump mstatus_csv_dumper_40;
    nodf_module_monitor module_monitor_40;
    nodf_module_intf module_intf_41(clock,reset);
    assign module_intf_41.ap_start = 1'b0;
    assign module_intf_41.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.tmp_47_modp_montymul_fu_3473.ap_ready;
    assign module_intf_41.ap_done = 1'b0;
    assign module_intf_41.ap_continue = 1'b0;
    assign module_intf_41.finish = finish;
    csv_file_dump mstatus_csv_dumper_41;
    nodf_module_monitor module_monitor_41;
    nodf_module_intf module_intf_42(clock,reset);
    assign module_intf_42.ap_start = 1'b0;
    assign module_intf_42.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.tmp_48_modp_montymul_fu_3482.ap_ready;
    assign module_intf_42.ap_done = 1'b0;
    assign module_intf_42.ap_continue = 1'b0;
    assign module_intf_42.finish = finish;
    csv_file_dump mstatus_csv_dumper_42;
    nodf_module_monitor module_monitor_42;
    nodf_module_intf module_intf_43(clock,reset);
    assign module_intf_43.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_start;
    assign module_intf_43.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ready;
    assign module_intf_43.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_done;
    assign module_intf_43.ap_continue = 1'b1;
    assign module_intf_43.finish = finish;
    csv_file_dump mstatus_csv_dumper_43;
    nodf_module_monitor module_monitor_43;
    nodf_module_intf module_intf_44(clock,reset);
    assign module_intf_44.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_fpr_of_fu_3517.ap_start;
    assign module_intf_44.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_fpr_of_fu_3517.ap_ready;
    assign module_intf_44.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_fpr_of_fu_3517.ap_done;
    assign module_intf_44.ap_continue = 1'b1;
    assign module_intf_44.finish = finish;
    csv_file_dump mstatus_csv_dumper_44;
    nodf_module_monitor module_monitor_44;
    nodf_module_intf module_intf_45(clock,reset);
    assign module_intf_45.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_start;
    assign module_intf_45.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ready;
    assign module_intf_45.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_done;
    assign module_intf_45.ap_continue = 1'b1;
    assign module_intf_45.finish = finish;
    csv_file_dump mstatus_csv_dumper_45;
    nodf_module_monitor module_monitor_45;
    nodf_module_intf module_intf_46(clock,reset);
    assign module_intf_46.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_fpr_rint_fu_3539.ap_start;
    assign module_intf_46.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_fpr_rint_fu_3539.ap_ready;
    assign module_intf_46.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_fpr_rint_fu_3539.ap_done;
    assign module_intf_46.ap_continue = 1'b1;
    assign module_intf_46.finish = finish;
    csv_file_dump mstatus_csv_dumper_46;
    nodf_module_monitor module_monitor_46;
    nodf_module_intf module_intf_47(clock,reset);
    assign module_intf_47.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_mod_small_signed_1_fu_3545.ap_start;
    assign module_intf_47.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_mod_small_signed_1_fu_3545.ap_ready;
    assign module_intf_47.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_mod_small_signed_1_fu_3545.ap_done;
    assign module_intf_47.ap_continue = 1'b1;
    assign module_intf_47.finish = finish;
    csv_file_dump mstatus_csv_dumper_47;
    nodf_module_monitor module_monitor_47;
    nodf_module_intf module_intf_48(clock,reset);
    assign module_intf_48.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_start;
    assign module_intf_48.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ready;
    assign module_intf_48.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_done;
    assign module_intf_48.ap_continue = 1'b1;
    assign module_intf_48.finish = finish;
    csv_file_dump mstatus_csv_dumper_48;
    nodf_module_monitor module_monitor_48;
    nodf_module_intf module_intf_49(clock,reset);
    assign module_intf_49.ap_start = 1'b0;
    assign module_intf_49.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.grp_modp_montymul_fu_442.ap_ready;
    assign module_intf_49.ap_done = 1'b0;
    assign module_intf_49.ap_continue = 1'b0;
    assign module_intf_49.finish = finish;
    csv_file_dump mstatus_csv_dumper_49;
    nodf_module_monitor module_monitor_49;
    nodf_module_intf module_intf_50(clock,reset);
    assign module_intf_50.ap_start = 1'b0;
    assign module_intf_50.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.grp_modp_montymul_fu_450.ap_ready;
    assign module_intf_50.ap_done = 1'b0;
    assign module_intf_50.ap_continue = 1'b0;
    assign module_intf_50.finish = finish;
    csv_file_dump mstatus_csv_dumper_50;
    nodf_module_monitor module_monitor_50;
    nodf_module_intf module_intf_51(clock,reset);
    assign module_intf_51.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_start;
    assign module_intf_51.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ready;
    assign module_intf_51.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_done;
    assign module_intf_51.ap_continue = 1'b1;
    assign module_intf_51.finish = finish;
    csv_file_dump mstatus_csv_dumper_51;
    nodf_module_monitor module_monitor_51;
    nodf_module_intf module_intf_52(clock,reset);
    assign module_intf_52.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.grp_fpr_of_fu_228.ap_start;
    assign module_intf_52.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.grp_fpr_of_fu_228.ap_ready;
    assign module_intf_52.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.grp_fpr_of_fu_228.ap_done;
    assign module_intf_52.ap_continue = 1'b1;
    assign module_intf_52.finish = finish;
    csv_file_dump mstatus_csv_dumper_52;
    nodf_module_monitor module_monitor_52;
    nodf_module_intf module_intf_53(clock,reset);
    assign module_intf_53.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_mul_fft_1_fu_3613.ap_start;
    assign module_intf_53.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_mul_fft_1_fu_3613.ap_ready;
    assign module_intf_53.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_mul_fft_1_fu_3613.ap_done;
    assign module_intf_53.ap_continue = 1'b1;
    assign module_intf_53.finish = finish;
    csv_file_dump mstatus_csv_dumper_53;
    nodf_module_monitor module_monitor_53;
    nodf_module_intf module_intf_54(clock,reset);
    assign module_intf_54.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_start;
    assign module_intf_54.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ready;
    assign module_intf_54.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_done;
    assign module_intf_54.ap_continue = 1'b1;
    assign module_intf_54.finish = finish;
    csv_file_dump mstatus_csv_dumper_54;
    nodf_module_monitor module_monitor_54;
    nodf_module_intf module_intf_55(clock,reset);
    assign module_intf_55.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_start;
    assign module_intf_55.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ready;
    assign module_intf_55.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_done;
    assign module_intf_55.ap_continue = 1'b1;
    assign module_intf_55.finish = finish;
    csv_file_dump mstatus_csv_dumper_55;
    nodf_module_monitor module_monitor_55;
    nodf_module_intf module_intf_56(clock,reset);
    assign module_intf_56.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_start;
    assign module_intf_56.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ready;
    assign module_intf_56.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_done;
    assign module_intf_56.ap_continue = 1'b1;
    assign module_intf_56.finish = finish;
    csv_file_dump mstatus_csv_dumper_56;
    nodf_module_monitor module_monitor_56;
    nodf_module_intf module_intf_57(clock,reset);
    assign module_intf_57.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_start;
    assign module_intf_57.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ready;
    assign module_intf_57.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_done;
    assign module_intf_57.ap_continue = 1'b1;
    assign module_intf_57.finish = finish;
    csv_file_dump mstatus_csv_dumper_57;
    nodf_module_monitor module_monitor_57;
    nodf_module_intf module_intf_58(clock,reset);
    assign module_intf_58.ap_start = 1'b0;
    assign module_intf_58.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_montymul_fu_800.ap_ready;
    assign module_intf_58.ap_done = 1'b0;
    assign module_intf_58.ap_continue = 1'b0;
    assign module_intf_58.finish = finish;
    csv_file_dump mstatus_csv_dumper_58;
    nodf_module_monitor module_monitor_58;
    nodf_module_intf module_intf_59(clock,reset);
    assign module_intf_59.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_start;
    assign module_intf_59.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ready;
    assign module_intf_59.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_done;
    assign module_intf_59.ap_continue = 1'b1;
    assign module_intf_59.finish = finish;
    csv_file_dump mstatus_csv_dumper_59;
    nodf_module_monitor module_monitor_59;
    nodf_module_intf module_intf_60(clock,reset);
    assign module_intf_60.ap_start = 1'b0;
    assign module_intf_60.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.grp_modp_montymul_fu_442.ap_ready;
    assign module_intf_60.ap_done = 1'b0;
    assign module_intf_60.ap_continue = 1'b0;
    assign module_intf_60.finish = finish;
    csv_file_dump mstatus_csv_dumper_60;
    nodf_module_monitor module_monitor_60;
    nodf_module_intf module_intf_61(clock,reset);
    assign module_intf_61.ap_start = 1'b0;
    assign module_intf_61.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.grp_modp_montymul_fu_450.ap_ready;
    assign module_intf_61.ap_done = 1'b0;
    assign module_intf_61.ap_continue = 1'b0;
    assign module_intf_61.finish = finish;
    csv_file_dump mstatus_csv_dumper_61;
    nodf_module_monitor module_monitor_61;
    nodf_module_intf module_intf_62(clock,reset);
    assign module_intf_62.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_start;
    assign module_intf_62.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ready;
    assign module_intf_62.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_done;
    assign module_intf_62.ap_continue = 1'b1;
    assign module_intf_62.finish = finish;
    csv_file_dump mstatus_csv_dumper_62;
    nodf_module_monitor module_monitor_62;
    nodf_module_intf module_intf_63(clock,reset);
    assign module_intf_63.ap_start = 1'b0;
    assign module_intf_63.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.y_modp_montymul_fu_200.ap_ready;
    assign module_intf_63.ap_done = 1'b0;
    assign module_intf_63.ap_continue = 1'b0;
    assign module_intf_63.finish = finish;
    csv_file_dump mstatus_csv_dumper_63;
    nodf_module_monitor module_monitor_63;
    nodf_module_intf module_intf_64(clock,reset);
    assign module_intf_64.ap_start = 1'b0;
    assign module_intf_64.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_montymul_fu_514.ap_ready;
    assign module_intf_64.ap_done = 1'b0;
    assign module_intf_64.ap_continue = 1'b0;
    assign module_intf_64.finish = finish;
    csv_file_dump mstatus_csv_dumper_64;
    nodf_module_monitor module_monitor_64;
    nodf_module_intf module_intf_65(clock,reset);
    assign module_intf_65.ap_start = 1'b0;
    assign module_intf_65.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_montymul_fu_524.ap_ready;
    assign module_intf_65.ap_done = 1'b0;
    assign module_intf_65.ap_continue = 1'b0;
    assign module_intf_65.finish = finish;
    csv_file_dump mstatus_csv_dumper_65;
    nodf_module_monitor module_monitor_65;
    nodf_module_intf module_intf_66(clock,reset);
    assign module_intf_66.ap_start = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_start;
    assign module_intf_66.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ready;
    assign module_intf_66.ap_done = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_done;
    assign module_intf_66.ap_continue = 1'b1;
    assign module_intf_66.finish = finish;
    csv_file_dump mstatus_csv_dumper_66;
    nodf_module_monitor module_monitor_66;
    nodf_module_intf module_intf_67(clock,reset);
    assign module_intf_67.ap_start = 1'b0;
    assign module_intf_67.ap_ready = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.y_modp_montymul_fu_200.ap_ready;
    assign module_intf_67.ap_done = 1'b0;
    assign module_intf_67.ap_continue = 1'b0;
    assign module_intf_67.finish = finish;
    csv_file_dump mstatus_csv_dumper_67;
    nodf_module_monitor module_monitor_67;

    seq_loop_intf#(117) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state1;
    assign seq_loop_intf_1.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_1.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state4;
    assign seq_loop_intf_1.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.post_loop_state1 = 117'h0;
    assign seq_loop_intf_1.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.post_loop_state2 = 117'h0;
    assign seq_loop_intf_1.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_1.post_loop_state3 = 117'h0;
    assign seq_loop_intf_1.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state2;
    assign seq_loop_intf_1.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_1.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state2;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state3;
    assign seq_loop_intf_1.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.iter_end_state1 = 117'h0;
    assign seq_loop_intf_1.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(117) seq_loop_monitor_1;
    seq_loop_intf#(117) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state2;
    assign seq_loop_intf_2.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_2.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state14;
    assign seq_loop_intf_2.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.post_loop_state1 = 117'h0;
    assign seq_loop_intf_2.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.post_loop_state2 = 117'h0;
    assign seq_loop_intf_2.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_2.post_loop_state3 = 117'h0;
    assign seq_loop_intf_2.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state4;
    assign seq_loop_intf_2.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_2.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state4;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state13;
    assign seq_loop_intf_2.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.iter_end_state1 = 117'h0;
    assign seq_loop_intf_2.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(117) seq_loop_monitor_2;
    seq_loop_intf#(117) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state16;
    assign seq_loop_intf_3.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_3.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state76;
    assign seq_loop_intf_3.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.post_loop_state1 = AESL_inst_keygen.ap_ST_fsm_state19;
    assign seq_loop_intf_3.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_3.post_loop_state2 = 117'h0;
    assign seq_loop_intf_3.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_3.post_loop_state3 = 117'h0;
    assign seq_loop_intf_3.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state17;
    assign seq_loop_intf_3.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_3.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state17;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state18;
    assign seq_loop_intf_3.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.iter_end_state1 = 117'h0;
    assign seq_loop_intf_3.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(117) seq_loop_monitor_3;
    seq_loop_intf#(117) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state17;
    assign seq_loop_intf_4.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_4.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state24;
    assign seq_loop_intf_4.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.post_loop_state1 = 117'h0;
    assign seq_loop_intf_4.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.post_loop_state2 = 117'h0;
    assign seq_loop_intf_4.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_4.post_loop_state3 = 117'h0;
    assign seq_loop_intf_4.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state19;
    assign seq_loop_intf_4.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_4.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state19;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state23;
    assign seq_loop_intf_4.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.iter_end_state1 = 117'h0;
    assign seq_loop_intf_4.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(117) seq_loop_monitor_4;
    seq_loop_intf#(117) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state19;
    assign seq_loop_intf_5.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_5.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state76;
    assign seq_loop_intf_5.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.post_loop_state1 = AESL_inst_keygen.ap_ST_fsm_state29;
    assign seq_loop_intf_5.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_5.post_loop_state2 = 117'h0;
    assign seq_loop_intf_5.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_5.post_loop_state3 = 117'h0;
    assign seq_loop_intf_5.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state24;
    assign seq_loop_intf_5.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_5.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state24;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state28;
    assign seq_loop_intf_5.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.iter_end_state1 = 117'h0;
    assign seq_loop_intf_5.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(117) seq_loop_monitor_5;
    seq_loop_intf#(117) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state24;
    assign seq_loop_intf_6.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_6.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state32;
    assign seq_loop_intf_6.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.post_loop_state1 = 117'h0;
    assign seq_loop_intf_6.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.post_loop_state2 = 117'h0;
    assign seq_loop_intf_6.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_6.post_loop_state3 = 117'h0;
    assign seq_loop_intf_6.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state29;
    assign seq_loop_intf_6.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_6.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state29;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state31;
    assign seq_loop_intf_6.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.iter_end_state1 = 117'h0;
    assign seq_loop_intf_6.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(117) seq_loop_monitor_6;
    seq_loop_intf#(117) seq_loop_intf_7(clock,reset);
    assign seq_loop_intf_7.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state29;
    assign seq_loop_intf_7.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_7.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state35;
    assign seq_loop_intf_7.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.post_loop_state1 = 117'h0;
    assign seq_loop_intf_7.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.post_loop_state2 = 117'h0;
    assign seq_loop_intf_7.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_7.post_loop_state3 = 117'h0;
    assign seq_loop_intf_7.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_7.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state32;
    assign seq_loop_intf_7.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_7.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_7.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state32;
    assign seq_loop_intf_7.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state34;
    assign seq_loop_intf_7.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.iter_end_state1 = 117'h0;
    assign seq_loop_intf_7.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.one_state_loop = 1'b0;
    assign seq_loop_intf_7.one_state_block = 1'b0;
    assign seq_loop_intf_7.finish = finish;
    csv_file_dump seq_loop_csv_dumper_7;
    seq_loop_monitor #(117) seq_loop_monitor_7;
    seq_loop_intf#(117) seq_loop_intf_8(clock,reset);
    assign seq_loop_intf_8.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state35;
    assign seq_loop_intf_8.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_8.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state48;
    assign seq_loop_intf_8.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.post_loop_state1 = 117'h0;
    assign seq_loop_intf_8.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.post_loop_state2 = 117'h0;
    assign seq_loop_intf_8.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_8.post_loop_state3 = 117'h0;
    assign seq_loop_intf_8.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_8.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state36;
    assign seq_loop_intf_8.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_8.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_8.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state36;
    assign seq_loop_intf_8.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state47;
    assign seq_loop_intf_8.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.iter_end_state1 = 117'h0;
    assign seq_loop_intf_8.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.one_state_loop = 1'b0;
    assign seq_loop_intf_8.one_state_block = 1'b0;
    assign seq_loop_intf_8.finish = finish;
    csv_file_dump seq_loop_csv_dumper_8;
    seq_loop_monitor #(117) seq_loop_monitor_8;
    seq_loop_intf#(117) seq_loop_intf_9(clock,reset);
    assign seq_loop_intf_9.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state36;
    assign seq_loop_intf_9.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_9.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state50;
    assign seq_loop_intf_9.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.post_loop_state1 = 117'h0;
    assign seq_loop_intf_9.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.post_loop_state2 = 117'h0;
    assign seq_loop_intf_9.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_9.post_loop_state3 = 117'h0;
    assign seq_loop_intf_9.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_9.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state48;
    assign seq_loop_intf_9.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_9.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_9.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state48;
    assign seq_loop_intf_9.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state49;
    assign seq_loop_intf_9.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.iter_end_state1 = 117'h0;
    assign seq_loop_intf_9.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.one_state_loop = 1'b0;
    assign seq_loop_intf_9.one_state_block = 1'b0;
    assign seq_loop_intf_9.finish = finish;
    csv_file_dump seq_loop_csv_dumper_9;
    seq_loop_monitor #(117) seq_loop_monitor_9;
    seq_loop_intf#(117) seq_loop_intf_10(clock,reset);
    assign seq_loop_intf_10.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state48;
    assign seq_loop_intf_10.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_10.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state52;
    assign seq_loop_intf_10.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.post_loop_state1 = 117'h0;
    assign seq_loop_intf_10.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.post_loop_state2 = 117'h0;
    assign seq_loop_intf_10.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_10.post_loop_state3 = 117'h0;
    assign seq_loop_intf_10.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_10.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state50;
    assign seq_loop_intf_10.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_10.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_10.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state50;
    assign seq_loop_intf_10.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state51;
    assign seq_loop_intf_10.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.iter_end_state1 = 117'h0;
    assign seq_loop_intf_10.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.one_state_loop = 1'b0;
    assign seq_loop_intf_10.one_state_block = 1'b0;
    assign seq_loop_intf_10.finish = finish;
    csv_file_dump seq_loop_csv_dumper_10;
    seq_loop_monitor #(117) seq_loop_monitor_10;
    seq_loop_intf#(117) seq_loop_intf_11(clock,reset);
    assign seq_loop_intf_11.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state50;
    assign seq_loop_intf_11.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_11.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state55;
    assign seq_loop_intf_11.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.post_loop_state1 = 117'h0;
    assign seq_loop_intf_11.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.post_loop_state2 = 117'h0;
    assign seq_loop_intf_11.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_11.post_loop_state3 = 117'h0;
    assign seq_loop_intf_11.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_11.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state52;
    assign seq_loop_intf_11.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_11.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_11.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state52;
    assign seq_loop_intf_11.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state54;
    assign seq_loop_intf_11.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.iter_end_state1 = 117'h0;
    assign seq_loop_intf_11.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.one_state_loop = 1'b0;
    assign seq_loop_intf_11.one_state_block = 1'b0;
    assign seq_loop_intf_11.finish = finish;
    csv_file_dump seq_loop_csv_dumper_11;
    seq_loop_monitor #(117) seq_loop_monitor_11;
    seq_loop_intf#(117) seq_loop_intf_12(clock,reset);
    assign seq_loop_intf_12.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state52;
    assign seq_loop_intf_12.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_12.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state58;
    assign seq_loop_intf_12.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.post_loop_state1 = 117'h0;
    assign seq_loop_intf_12.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.post_loop_state2 = 117'h0;
    assign seq_loop_intf_12.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_12.post_loop_state3 = 117'h0;
    assign seq_loop_intf_12.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_12.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state55;
    assign seq_loop_intf_12.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_12.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_12.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state55;
    assign seq_loop_intf_12.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state57;
    assign seq_loop_intf_12.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.iter_end_state1 = 117'h0;
    assign seq_loop_intf_12.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.one_state_loop = 1'b0;
    assign seq_loop_intf_12.one_state_block = 1'b0;
    assign seq_loop_intf_12.finish = finish;
    csv_file_dump seq_loop_csv_dumper_12;
    seq_loop_monitor #(117) seq_loop_monitor_12;
    seq_loop_intf#(117) seq_loop_intf_13(clock,reset);
    assign seq_loop_intf_13.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state55;
    assign seq_loop_intf_13.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_13.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state61;
    assign seq_loop_intf_13.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.post_loop_state1 = 117'h0;
    assign seq_loop_intf_13.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.post_loop_state2 = 117'h0;
    assign seq_loop_intf_13.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_13.post_loop_state3 = 117'h0;
    assign seq_loop_intf_13.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_13.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state58;
    assign seq_loop_intf_13.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_13.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_13.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state58;
    assign seq_loop_intf_13.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state60;
    assign seq_loop_intf_13.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.iter_end_state1 = 117'h0;
    assign seq_loop_intf_13.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.one_state_loop = 1'b0;
    assign seq_loop_intf_13.one_state_block = 1'b0;
    assign seq_loop_intf_13.finish = finish;
    csv_file_dump seq_loop_csv_dumper_13;
    seq_loop_monitor #(117) seq_loop_monitor_13;
    seq_loop_intf#(117) seq_loop_intf_14(clock,reset);
    assign seq_loop_intf_14.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state58;
    assign seq_loop_intf_14.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_14.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state64;
    assign seq_loop_intf_14.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.post_loop_state1 = 117'h0;
    assign seq_loop_intf_14.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.post_loop_state2 = 117'h0;
    assign seq_loop_intf_14.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_14.post_loop_state3 = 117'h0;
    assign seq_loop_intf_14.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_14.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state61;
    assign seq_loop_intf_14.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_14.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_14.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state61;
    assign seq_loop_intf_14.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state63;
    assign seq_loop_intf_14.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.iter_end_state1 = 117'h0;
    assign seq_loop_intf_14.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_14.one_state_loop = 1'b0;
    assign seq_loop_intf_14.one_state_block = 1'b0;
    assign seq_loop_intf_14.finish = finish;
    csv_file_dump seq_loop_csv_dumper_14;
    seq_loop_monitor #(117) seq_loop_monitor_14;
    seq_loop_intf#(117) seq_loop_intf_15(clock,reset);
    assign seq_loop_intf_15.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state64;
    assign seq_loop_intf_15.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_15.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state71;
    assign seq_loop_intf_15.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.post_loop_state1 = 117'h0;
    assign seq_loop_intf_15.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.post_loop_state2 = 117'h0;
    assign seq_loop_intf_15.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_15.post_loop_state3 = 117'h0;
    assign seq_loop_intf_15.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_15.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state65;
    assign seq_loop_intf_15.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_15.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_15.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state65;
    assign seq_loop_intf_15.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state70;
    assign seq_loop_intf_15.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.iter_end_state1 = 117'h0;
    assign seq_loop_intf_15.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.one_state_loop = 1'b0;
    assign seq_loop_intf_15.one_state_block = 1'b0;
    assign seq_loop_intf_15.finish = finish;
    csv_file_dump seq_loop_csv_dumper_15;
    seq_loop_monitor #(117) seq_loop_monitor_15;
    seq_loop_intf#(117) seq_loop_intf_16(clock,reset);
    assign seq_loop_intf_16.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state4;
    assign seq_loop_intf_16.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_16.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_16.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state77;
    assign seq_loop_intf_16.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.post_loop_state1 = 117'h0;
    assign seq_loop_intf_16.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_16.post_loop_state2 = 117'h0;
    assign seq_loop_intf_16.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_16.post_loop_state3 = 117'h0;
    assign seq_loop_intf_16.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_16.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state76;
    assign seq_loop_intf_16.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_16.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_16.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_16.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state14;
    assign seq_loop_intf_16.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state76;
    assign seq_loop_intf_16.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.iter_end_state1 = 117'h0;
    assign seq_loop_intf_16.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_16.one_state_loop = 1'b0;
    assign seq_loop_intf_16.one_state_block = 1'b0;
    assign seq_loop_intf_16.finish = finish;
    csv_file_dump seq_loop_csv_dumper_16;
    seq_loop_monitor #(117) seq_loop_monitor_16;
    seq_loop_intf#(117) seq_loop_intf_17(clock,reset);
    assign seq_loop_intf_17.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state76;
    assign seq_loop_intf_17.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_17.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_17.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state85;
    assign seq_loop_intf_17.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.post_loop_state1 = 117'h0;
    assign seq_loop_intf_17.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_17.post_loop_state2 = 117'h0;
    assign seq_loop_intf_17.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_17.post_loop_state3 = 117'h0;
    assign seq_loop_intf_17.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_17.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state77;
    assign seq_loop_intf_17.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_17.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_17.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_17.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state77;
    assign seq_loop_intf_17.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state84;
    assign seq_loop_intf_17.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.iter_end_state1 = 117'h0;
    assign seq_loop_intf_17.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_17.one_state_loop = 1'b0;
    assign seq_loop_intf_17.one_state_block = 1'b0;
    assign seq_loop_intf_17.finish = finish;
    csv_file_dump seq_loop_csv_dumper_17;
    seq_loop_monitor #(117) seq_loop_monitor_17;
    seq_loop_intf#(117) seq_loop_intf_18(clock,reset);
    assign seq_loop_intf_18.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state77;
    assign seq_loop_intf_18.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_18.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_18.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_18.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state93;
    assign seq_loop_intf_18.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_18.post_loop_state1 = 117'h0;
    assign seq_loop_intf_18.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_18.post_loop_state2 = 117'h0;
    assign seq_loop_intf_18.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_18.post_loop_state3 = 117'h0;
    assign seq_loop_intf_18.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_18.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state85;
    assign seq_loop_intf_18.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_18.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_18.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_18.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_18.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state85;
    assign seq_loop_intf_18.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state92;
    assign seq_loop_intf_18.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_18.iter_end_state1 = 117'h0;
    assign seq_loop_intf_18.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_18.one_state_loop = 1'b0;
    assign seq_loop_intf_18.one_state_block = 1'b0;
    assign seq_loop_intf_18.finish = finish;
    csv_file_dump seq_loop_csv_dumper_18;
    seq_loop_monitor #(117) seq_loop_monitor_18;
    seq_loop_intf#(117) seq_loop_intf_19(clock,reset);
    assign seq_loop_intf_19.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state93;
    assign seq_loop_intf_19.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_19.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_19.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_19.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state97;
    assign seq_loop_intf_19.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_19.post_loop_state1 = 117'h0;
    assign seq_loop_intf_19.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_19.post_loop_state2 = 117'h0;
    assign seq_loop_intf_19.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_19.post_loop_state3 = 117'h0;
    assign seq_loop_intf_19.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_19.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state94;
    assign seq_loop_intf_19.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_19.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_19.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_19.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_19.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state94;
    assign seq_loop_intf_19.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state96;
    assign seq_loop_intf_19.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_19.iter_end_state1 = 117'h0;
    assign seq_loop_intf_19.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_19.one_state_loop = 1'b0;
    assign seq_loop_intf_19.one_state_block = 1'b0;
    assign seq_loop_intf_19.finish = finish;
    csv_file_dump seq_loop_csv_dumper_19;
    seq_loop_monitor #(117) seq_loop_monitor_19;
    seq_loop_intf#(117) seq_loop_intf_20(clock,reset);
    assign seq_loop_intf_20.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state101;
    assign seq_loop_intf_20.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_20.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_20.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_20.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state110;
    assign seq_loop_intf_20.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_20.post_loop_state1 = 117'h0;
    assign seq_loop_intf_20.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_20.post_loop_state2 = 117'h0;
    assign seq_loop_intf_20.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_20.post_loop_state3 = 117'h0;
    assign seq_loop_intf_20.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_20.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state102;
    assign seq_loop_intf_20.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_20.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_20.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_20.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_20.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state102;
    assign seq_loop_intf_20.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state109;
    assign seq_loop_intf_20.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_20.iter_end_state1 = 117'h0;
    assign seq_loop_intf_20.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_20.one_state_loop = 1'b0;
    assign seq_loop_intf_20.one_state_block = 1'b0;
    assign seq_loop_intf_20.finish = finish;
    csv_file_dump seq_loop_csv_dumper_20;
    seq_loop_monitor #(117) seq_loop_monitor_20;
    seq_loop_intf#(117) seq_loop_intf_21(clock,reset);
    assign seq_loop_intf_21.pre_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state102;
    assign seq_loop_intf_21.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_21.pre_loop_state1 = 117'h0;
    assign seq_loop_intf_21.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_21.post_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state1;
    assign seq_loop_intf_21.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_21.post_loop_state1 = 117'h0;
    assign seq_loop_intf_21.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_21.post_loop_state2 = 117'h0;
    assign seq_loop_intf_21.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_21.post_loop_state3 = 117'h0;
    assign seq_loop_intf_21.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_21.quit_loop_state0 = AESL_inst_keygen.ap_ST_fsm_state110;
    assign seq_loop_intf_21.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_21.quit_loop_state1 = 117'h0;
    assign seq_loop_intf_21.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_21.cur_state = AESL_inst_keygen.ap_CS_fsm;
    assign seq_loop_intf_21.iter_start_state = AESL_inst_keygen.ap_ST_fsm_state110;
    assign seq_loop_intf_21.iter_end_state0 = AESL_inst_keygen.ap_ST_fsm_state117;
    assign seq_loop_intf_21.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_21.iter_end_state1 = 117'h0;
    assign seq_loop_intf_21.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_21.one_state_loop = 1'b0;
    assign seq_loop_intf_21.one_state_block = 1'b0;
    assign seq_loop_intf_21.finish = finish;
    csv_file_dump seq_loop_csv_dumper_21;
    seq_loop_monitor #(117) seq_loop_monitor_21;
    seq_loop_intf#(7) seq_loop_intf_22(clock,reset);
    assign seq_loop_intf_22.pre_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state5;
    assign seq_loop_intf_22.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_22.pre_loop_state1 = 7'h0;
    assign seq_loop_intf_22.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_22.post_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state2;
    assign seq_loop_intf_22.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_22.post_loop_state1 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state3;
    assign seq_loop_intf_22.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_22.post_loop_state2 = 7'h0;
    assign seq_loop_intf_22.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_22.post_loop_state3 = 7'h0;
    assign seq_loop_intf_22.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_22.quit_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state6;
    assign seq_loop_intf_22.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_22.quit_loop_state1 = 7'h0;
    assign seq_loop_intf_22.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_22.cur_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_CS_fsm;
    assign seq_loop_intf_22.iter_start_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state6;
    assign seq_loop_intf_22.iter_end_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state7;
    assign seq_loop_intf_22.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_22.iter_end_state1 = 7'h0;
    assign seq_loop_intf_22.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_22.one_state_loop = 1'b0;
    assign seq_loop_intf_22.one_state_block = 1'b0;
    assign seq_loop_intf_22.finish = finish;
    csv_file_dump seq_loop_csv_dumper_22;
    seq_loop_monitor #(7) seq_loop_monitor_22;
    seq_loop_intf#(7) seq_loop_intf_23(clock,reset);
    assign seq_loop_intf_23.pre_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state2;
    assign seq_loop_intf_23.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_23.pre_loop_state1 = 7'h0;
    assign seq_loop_intf_23.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_23.post_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state2;
    assign seq_loop_intf_23.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_23.post_loop_state1 = 7'h0;
    assign seq_loop_intf_23.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_23.post_loop_state2 = 7'h0;
    assign seq_loop_intf_23.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_23.post_loop_state3 = 7'h0;
    assign seq_loop_intf_23.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_23.quit_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state6;
    assign seq_loop_intf_23.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_23.quit_loop_state1 = 7'h0;
    assign seq_loop_intf_23.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_23.cur_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_CS_fsm;
    assign seq_loop_intf_23.iter_start_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state3;
    assign seq_loop_intf_23.iter_end_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state6;
    assign seq_loop_intf_23.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_23.iter_end_state1 = 7'h0;
    assign seq_loop_intf_23.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_23.one_state_loop = 1'b0;
    assign seq_loop_intf_23.one_state_block = 1'b0;
    assign seq_loop_intf_23.finish = finish;
    csv_file_dump seq_loop_csv_dumper_23;
    seq_loop_monitor #(7) seq_loop_monitor_23;
    seq_loop_intf#(7) seq_loop_intf_24(clock,reset);
    assign seq_loop_intf_24.pre_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state1;
    assign seq_loop_intf_24.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_24.pre_loop_state1 = 7'h0;
    assign seq_loop_intf_24.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_24.post_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state1;
    assign seq_loop_intf_24.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_24.post_loop_state1 = 7'h0;
    assign seq_loop_intf_24.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_24.post_loop_state2 = 7'h0;
    assign seq_loop_intf_24.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_24.post_loop_state3 = 7'h0;
    assign seq_loop_intf_24.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_24.quit_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state2;
    assign seq_loop_intf_24.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_24.quit_loop_state1 = 7'h0;
    assign seq_loop_intf_24.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_24.cur_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_CS_fsm;
    assign seq_loop_intf_24.iter_start_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state2;
    assign seq_loop_intf_24.iter_end_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.ap_ST_fsm_state6;
    assign seq_loop_intf_24.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_24.iter_end_state1 = 7'h0;
    assign seq_loop_intf_24.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_24.one_state_loop = 1'b0;
    assign seq_loop_intf_24.one_state_block = 1'b0;
    assign seq_loop_intf_24.finish = finish;
    csv_file_dump seq_loop_csv_dumper_24;
    seq_loop_monitor #(7) seq_loop_monitor_24;
    seq_loop_intf#(10) seq_loop_intf_25(clock,reset);
    assign seq_loop_intf_25.pre_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state4;
    assign seq_loop_intf_25.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_25.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_25.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_25.post_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state6;
    assign seq_loop_intf_25.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_25.post_loop_state1 = 10'h0;
    assign seq_loop_intf_25.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_25.post_loop_state2 = 10'h0;
    assign seq_loop_intf_25.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_25.post_loop_state3 = 10'h0;
    assign seq_loop_intf_25.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_25.quit_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state5;
    assign seq_loop_intf_25.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_25.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_25.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_25.cur_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_CS_fsm;
    assign seq_loop_intf_25.iter_start_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state5;
    assign seq_loop_intf_25.iter_end_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state5;
    assign seq_loop_intf_25.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_25.iter_end_state1 = 10'h0;
    assign seq_loop_intf_25.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_25.one_state_loop = 1'b1;
    assign seq_loop_intf_25.one_state_block = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state5_blk;
    assign seq_loop_intf_25.finish = finish;
    csv_file_dump seq_loop_csv_dumper_25;
    seq_loop_monitor #(10) seq_loop_monitor_25;
    seq_loop_intf#(10) seq_loop_intf_26(clock,reset);
    assign seq_loop_intf_26.pre_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state1;
    assign seq_loop_intf_26.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_26.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_26.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_26.post_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state7;
    assign seq_loop_intf_26.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_26.post_loop_state1 = 10'h0;
    assign seq_loop_intf_26.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_26.post_loop_state2 = 10'h0;
    assign seq_loop_intf_26.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_26.post_loop_state3 = 10'h0;
    assign seq_loop_intf_26.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_26.quit_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state2;
    assign seq_loop_intf_26.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_26.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_26.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_26.cur_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_CS_fsm;
    assign seq_loop_intf_26.iter_start_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state2;
    assign seq_loop_intf_26.iter_end_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.ap_ST_fsm_state6;
    assign seq_loop_intf_26.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_26.iter_end_state1 = 10'h0;
    assign seq_loop_intf_26.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_26.one_state_loop = 1'b0;
    assign seq_loop_intf_26.one_state_block = 1'b0;
    assign seq_loop_intf_26.finish = finish;
    csv_file_dump seq_loop_csv_dumper_26;
    seq_loop_monitor #(10) seq_loop_monitor_26;
    seq_loop_intf#(3) seq_loop_intf_27(clock,reset);
    assign seq_loop_intf_27.pre_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.grp_process_block_111_112_fu_512.ap_ST_fsm_state1;
    assign seq_loop_intf_27.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_27.pre_loop_state1 = 3'h0;
    assign seq_loop_intf_27.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_27.post_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.grp_process_block_111_112_fu_512.ap_ST_fsm_state1;
    assign seq_loop_intf_27.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_27.post_loop_state1 = 3'h0;
    assign seq_loop_intf_27.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_27.post_loop_state2 = 3'h0;
    assign seq_loop_intf_27.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_27.post_loop_state3 = 3'h0;
    assign seq_loop_intf_27.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_27.quit_loop_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.grp_process_block_111_112_fu_512.ap_ST_fsm_state2;
    assign seq_loop_intf_27.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_27.quit_loop_state1 = 3'h0;
    assign seq_loop_intf_27.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_27.cur_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.grp_process_block_111_112_fu_512.ap_CS_fsm;
    assign seq_loop_intf_27.iter_start_state = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.grp_process_block_111_112_fu_512.ap_ST_fsm_state2;
    assign seq_loop_intf_27.iter_end_state0 = AESL_inst_keygen.grp_poly_small_mkgauss_fu_1282.grp_get_rng_u64_82_101_fu_718.grp_process_block_111_112_fu_512.ap_ST_fsm_state3;
    assign seq_loop_intf_27.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_27.iter_end_state1 = 3'h0;
    assign seq_loop_intf_27.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_27.one_state_loop = 1'b0;
    assign seq_loop_intf_27.one_state_block = 1'b0;
    assign seq_loop_intf_27.finish = finish;
    csv_file_dump seq_loop_csv_dumper_27;
    seq_loop_monitor #(3) seq_loop_monitor_27;
    seq_loop_intf#(10) seq_loop_intf_28(clock,reset);
    assign seq_loop_intf_28.pre_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state4;
    assign seq_loop_intf_28.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_28.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_28.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_28.post_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state3;
    assign seq_loop_intf_28.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_28.post_loop_state1 = 10'h0;
    assign seq_loop_intf_28.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_28.post_loop_state2 = 10'h0;
    assign seq_loop_intf_28.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_28.post_loop_state3 = 10'h0;
    assign seq_loop_intf_28.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_28.quit_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state5;
    assign seq_loop_intf_28.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_28.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_28.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_28.cur_state = AESL_inst_keygen.grp_FFT_fu_1324.ap_CS_fsm;
    assign seq_loop_intf_28.iter_start_state = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state5;
    assign seq_loop_intf_28.iter_end_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state10;
    assign seq_loop_intf_28.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_28.iter_end_state1 = 10'h0;
    assign seq_loop_intf_28.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_28.one_state_loop = 1'b0;
    assign seq_loop_intf_28.one_state_block = 1'b0;
    assign seq_loop_intf_28.finish = finish;
    csv_file_dump seq_loop_csv_dumper_28;
    seq_loop_monitor #(10) seq_loop_monitor_28;
    seq_loop_intf#(10) seq_loop_intf_29(clock,reset);
    assign seq_loop_intf_29.pre_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state2;
    assign seq_loop_intf_29.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_29.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_29.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_29.post_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state2;
    assign seq_loop_intf_29.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_29.post_loop_state1 = 10'h0;
    assign seq_loop_intf_29.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_29.post_loop_state2 = 10'h0;
    assign seq_loop_intf_29.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_29.post_loop_state3 = 10'h0;
    assign seq_loop_intf_29.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_29.quit_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state3;
    assign seq_loop_intf_29.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_29.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_29.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_29.cur_state = AESL_inst_keygen.grp_FFT_fu_1324.ap_CS_fsm;
    assign seq_loop_intf_29.iter_start_state = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state3;
    assign seq_loop_intf_29.iter_end_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state5;
    assign seq_loop_intf_29.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_29.iter_end_state1 = 10'h0;
    assign seq_loop_intf_29.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_29.one_state_loop = 1'b0;
    assign seq_loop_intf_29.one_state_block = 1'b0;
    assign seq_loop_intf_29.finish = finish;
    csv_file_dump seq_loop_csv_dumper_29;
    seq_loop_monitor #(10) seq_loop_monitor_29;
    seq_loop_intf#(10) seq_loop_intf_30(clock,reset);
    assign seq_loop_intf_30.pre_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state1;
    assign seq_loop_intf_30.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_30.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_30.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_30.post_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state1;
    assign seq_loop_intf_30.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_30.post_loop_state1 = 10'h0;
    assign seq_loop_intf_30.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_30.post_loop_state2 = 10'h0;
    assign seq_loop_intf_30.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_30.post_loop_state3 = 10'h0;
    assign seq_loop_intf_30.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_30.quit_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state2;
    assign seq_loop_intf_30.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_30.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_30.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_30.cur_state = AESL_inst_keygen.grp_FFT_fu_1324.ap_CS_fsm;
    assign seq_loop_intf_30.iter_start_state = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state2;
    assign seq_loop_intf_30.iter_end_state0 = AESL_inst_keygen.grp_FFT_fu_1324.ap_ST_fsm_state3;
    assign seq_loop_intf_30.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_30.iter_end_state1 = 10'h0;
    assign seq_loop_intf_30.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_30.one_state_loop = 1'b0;
    assign seq_loop_intf_30.one_state_block = 1'b0;
    assign seq_loop_intf_30.finish = finish;
    csv_file_dump seq_loop_csv_dumper_30;
    seq_loop_monitor #(10) seq_loop_monitor_30;
    seq_loop_intf#(10) seq_loop_intf_31(clock,reset);
    assign seq_loop_intf_31.pre_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state4;
    assign seq_loop_intf_31.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_31.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_31.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_31.post_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state3;
    assign seq_loop_intf_31.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_31.post_loop_state1 = 10'h0;
    assign seq_loop_intf_31.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_31.post_loop_state2 = 10'h0;
    assign seq_loop_intf_31.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_31.post_loop_state3 = 10'h0;
    assign seq_loop_intf_31.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_31.quit_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state5;
    assign seq_loop_intf_31.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_31.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_31.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_31.cur_state = AESL_inst_keygen.grp_FFT_fu_1331.ap_CS_fsm;
    assign seq_loop_intf_31.iter_start_state = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state5;
    assign seq_loop_intf_31.iter_end_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state10;
    assign seq_loop_intf_31.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_31.iter_end_state1 = 10'h0;
    assign seq_loop_intf_31.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_31.one_state_loop = 1'b0;
    assign seq_loop_intf_31.one_state_block = 1'b0;
    assign seq_loop_intf_31.finish = finish;
    csv_file_dump seq_loop_csv_dumper_31;
    seq_loop_monitor #(10) seq_loop_monitor_31;
    seq_loop_intf#(10) seq_loop_intf_32(clock,reset);
    assign seq_loop_intf_32.pre_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state2;
    assign seq_loop_intf_32.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_32.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_32.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_32.post_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state2;
    assign seq_loop_intf_32.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_32.post_loop_state1 = 10'h0;
    assign seq_loop_intf_32.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_32.post_loop_state2 = 10'h0;
    assign seq_loop_intf_32.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_32.post_loop_state3 = 10'h0;
    assign seq_loop_intf_32.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_32.quit_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state3;
    assign seq_loop_intf_32.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_32.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_32.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_32.cur_state = AESL_inst_keygen.grp_FFT_fu_1331.ap_CS_fsm;
    assign seq_loop_intf_32.iter_start_state = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state3;
    assign seq_loop_intf_32.iter_end_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state5;
    assign seq_loop_intf_32.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_32.iter_end_state1 = 10'h0;
    assign seq_loop_intf_32.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_32.one_state_loop = 1'b0;
    assign seq_loop_intf_32.one_state_block = 1'b0;
    assign seq_loop_intf_32.finish = finish;
    csv_file_dump seq_loop_csv_dumper_32;
    seq_loop_monitor #(10) seq_loop_monitor_32;
    seq_loop_intf#(10) seq_loop_intf_33(clock,reset);
    assign seq_loop_intf_33.pre_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state1;
    assign seq_loop_intf_33.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_33.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_33.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_33.post_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state1;
    assign seq_loop_intf_33.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_33.post_loop_state1 = 10'h0;
    assign seq_loop_intf_33.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_33.post_loop_state2 = 10'h0;
    assign seq_loop_intf_33.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_33.post_loop_state3 = 10'h0;
    assign seq_loop_intf_33.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_33.quit_loop_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state2;
    assign seq_loop_intf_33.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_33.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_33.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_33.cur_state = AESL_inst_keygen.grp_FFT_fu_1331.ap_CS_fsm;
    assign seq_loop_intf_33.iter_start_state = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state2;
    assign seq_loop_intf_33.iter_end_state0 = AESL_inst_keygen.grp_FFT_fu_1331.ap_ST_fsm_state3;
    assign seq_loop_intf_33.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_33.iter_end_state1 = 10'h0;
    assign seq_loop_intf_33.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_33.one_state_loop = 1'b0;
    assign seq_loop_intf_33.one_state_block = 1'b0;
    assign seq_loop_intf_33.finish = finish;
    csv_file_dump seq_loop_csv_dumper_33;
    seq_loop_monitor #(10) seq_loop_monitor_33;
    seq_loop_intf#(13) seq_loop_intf_34(clock,reset);
    assign seq_loop_intf_34.pre_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state4;
    assign seq_loop_intf_34.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_34.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_34.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_34.post_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state3;
    assign seq_loop_intf_34.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_34.post_loop_state1 = 13'h0;
    assign seq_loop_intf_34.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_34.post_loop_state2 = 13'h0;
    assign seq_loop_intf_34.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_34.post_loop_state3 = 13'h0;
    assign seq_loop_intf_34.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_34.quit_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state5;
    assign seq_loop_intf_34.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_34.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_34.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_34.cur_state = AESL_inst_keygen.grp_iFFT_fu_1338.ap_CS_fsm;
    assign seq_loop_intf_34.iter_start_state = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state5;
    assign seq_loop_intf_34.iter_end_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state10;
    assign seq_loop_intf_34.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_34.iter_end_state1 = 13'h0;
    assign seq_loop_intf_34.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_34.one_state_loop = 1'b0;
    assign seq_loop_intf_34.one_state_block = 1'b0;
    assign seq_loop_intf_34.finish = finish;
    csv_file_dump seq_loop_csv_dumper_34;
    seq_loop_monitor #(13) seq_loop_monitor_34;
    seq_loop_intf#(13) seq_loop_intf_35(clock,reset);
    assign seq_loop_intf_35.pre_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state2;
    assign seq_loop_intf_35.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_35.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_35.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_35.post_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state2;
    assign seq_loop_intf_35.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_35.post_loop_state1 = 13'h0;
    assign seq_loop_intf_35.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_35.post_loop_state2 = 13'h0;
    assign seq_loop_intf_35.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_35.post_loop_state3 = 13'h0;
    assign seq_loop_intf_35.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_35.quit_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state3;
    assign seq_loop_intf_35.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_35.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_35.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_35.cur_state = AESL_inst_keygen.grp_iFFT_fu_1338.ap_CS_fsm;
    assign seq_loop_intf_35.iter_start_state = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state3;
    assign seq_loop_intf_35.iter_end_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state5;
    assign seq_loop_intf_35.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_35.iter_end_state1 = 13'h0;
    assign seq_loop_intf_35.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_35.one_state_loop = 1'b0;
    assign seq_loop_intf_35.one_state_block = 1'b0;
    assign seq_loop_intf_35.finish = finish;
    csv_file_dump seq_loop_csv_dumper_35;
    seq_loop_monitor #(13) seq_loop_monitor_35;
    seq_loop_intf#(13) seq_loop_intf_36(clock,reset);
    assign seq_loop_intf_36.pre_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state1;
    assign seq_loop_intf_36.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_36.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_36.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_36.post_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state11;
    assign seq_loop_intf_36.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_36.post_loop_state1 = 13'h0;
    assign seq_loop_intf_36.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_36.post_loop_state2 = 13'h0;
    assign seq_loop_intf_36.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_36.post_loop_state3 = 13'h0;
    assign seq_loop_intf_36.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_36.quit_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state2;
    assign seq_loop_intf_36.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_36.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_36.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_36.cur_state = AESL_inst_keygen.grp_iFFT_fu_1338.ap_CS_fsm;
    assign seq_loop_intf_36.iter_start_state = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state2;
    assign seq_loop_intf_36.iter_end_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state3;
    assign seq_loop_intf_36.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_36.iter_end_state1 = 13'h0;
    assign seq_loop_intf_36.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_36.one_state_loop = 1'b0;
    assign seq_loop_intf_36.one_state_block = 1'b0;
    assign seq_loop_intf_36.finish = finish;
    csv_file_dump seq_loop_csv_dumper_36;
    seq_loop_monitor #(13) seq_loop_monitor_36;
    seq_loop_intf#(13) seq_loop_intf_37(clock,reset);
    assign seq_loop_intf_37.pre_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state2;
    assign seq_loop_intf_37.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_37.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_37.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_37.post_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state1;
    assign seq_loop_intf_37.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_37.post_loop_state1 = 13'h0;
    assign seq_loop_intf_37.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_37.post_loop_state2 = 13'h0;
    assign seq_loop_intf_37.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_37.post_loop_state3 = 13'h0;
    assign seq_loop_intf_37.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_37.quit_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state11;
    assign seq_loop_intf_37.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_37.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_37.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_37.cur_state = AESL_inst_keygen.grp_iFFT_fu_1338.ap_CS_fsm;
    assign seq_loop_intf_37.iter_start_state = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state11;
    assign seq_loop_intf_37.iter_end_state0 = AESL_inst_keygen.grp_iFFT_fu_1338.ap_ST_fsm_state13;
    assign seq_loop_intf_37.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_37.iter_end_state1 = 13'h0;
    assign seq_loop_intf_37.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_37.one_state_loop = 1'b0;
    assign seq_loop_intf_37.one_state_block = 1'b0;
    assign seq_loop_intf_37.finish = finish;
    csv_file_dump seq_loop_csv_dumper_37;
    seq_loop_monitor #(13) seq_loop_monitor_37;
    seq_loop_intf#(13) seq_loop_intf_38(clock,reset);
    assign seq_loop_intf_38.pre_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state4;
    assign seq_loop_intf_38.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_38.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_38.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_38.post_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state3;
    assign seq_loop_intf_38.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_38.post_loop_state1 = 13'h0;
    assign seq_loop_intf_38.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_38.post_loop_state2 = 13'h0;
    assign seq_loop_intf_38.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_38.post_loop_state3 = 13'h0;
    assign seq_loop_intf_38.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_38.quit_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state5;
    assign seq_loop_intf_38.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_38.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_38.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_38.cur_state = AESL_inst_keygen.grp_iFFT_fu_1345.ap_CS_fsm;
    assign seq_loop_intf_38.iter_start_state = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state5;
    assign seq_loop_intf_38.iter_end_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state10;
    assign seq_loop_intf_38.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_38.iter_end_state1 = 13'h0;
    assign seq_loop_intf_38.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_38.one_state_loop = 1'b0;
    assign seq_loop_intf_38.one_state_block = 1'b0;
    assign seq_loop_intf_38.finish = finish;
    csv_file_dump seq_loop_csv_dumper_38;
    seq_loop_monitor #(13) seq_loop_monitor_38;
    seq_loop_intf#(13) seq_loop_intf_39(clock,reset);
    assign seq_loop_intf_39.pre_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state2;
    assign seq_loop_intf_39.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_39.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_39.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_39.post_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state2;
    assign seq_loop_intf_39.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_39.post_loop_state1 = 13'h0;
    assign seq_loop_intf_39.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_39.post_loop_state2 = 13'h0;
    assign seq_loop_intf_39.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_39.post_loop_state3 = 13'h0;
    assign seq_loop_intf_39.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_39.quit_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state3;
    assign seq_loop_intf_39.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_39.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_39.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_39.cur_state = AESL_inst_keygen.grp_iFFT_fu_1345.ap_CS_fsm;
    assign seq_loop_intf_39.iter_start_state = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state3;
    assign seq_loop_intf_39.iter_end_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state5;
    assign seq_loop_intf_39.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_39.iter_end_state1 = 13'h0;
    assign seq_loop_intf_39.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_39.one_state_loop = 1'b0;
    assign seq_loop_intf_39.one_state_block = 1'b0;
    assign seq_loop_intf_39.finish = finish;
    csv_file_dump seq_loop_csv_dumper_39;
    seq_loop_monitor #(13) seq_loop_monitor_39;
    seq_loop_intf#(13) seq_loop_intf_40(clock,reset);
    assign seq_loop_intf_40.pre_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state1;
    assign seq_loop_intf_40.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_40.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_40.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_40.post_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state11;
    assign seq_loop_intf_40.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_40.post_loop_state1 = 13'h0;
    assign seq_loop_intf_40.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_40.post_loop_state2 = 13'h0;
    assign seq_loop_intf_40.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_40.post_loop_state3 = 13'h0;
    assign seq_loop_intf_40.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_40.quit_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state2;
    assign seq_loop_intf_40.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_40.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_40.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_40.cur_state = AESL_inst_keygen.grp_iFFT_fu_1345.ap_CS_fsm;
    assign seq_loop_intf_40.iter_start_state = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state2;
    assign seq_loop_intf_40.iter_end_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state3;
    assign seq_loop_intf_40.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_40.iter_end_state1 = 13'h0;
    assign seq_loop_intf_40.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_40.one_state_loop = 1'b0;
    assign seq_loop_intf_40.one_state_block = 1'b0;
    assign seq_loop_intf_40.finish = finish;
    csv_file_dump seq_loop_csv_dumper_40;
    seq_loop_monitor #(13) seq_loop_monitor_40;
    seq_loop_intf#(13) seq_loop_intf_41(clock,reset);
    assign seq_loop_intf_41.pre_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state2;
    assign seq_loop_intf_41.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_41.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_41.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_41.post_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state1;
    assign seq_loop_intf_41.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_41.post_loop_state1 = 13'h0;
    assign seq_loop_intf_41.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_41.post_loop_state2 = 13'h0;
    assign seq_loop_intf_41.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_41.post_loop_state3 = 13'h0;
    assign seq_loop_intf_41.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_41.quit_loop_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state11;
    assign seq_loop_intf_41.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_41.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_41.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_41.cur_state = AESL_inst_keygen.grp_iFFT_fu_1345.ap_CS_fsm;
    assign seq_loop_intf_41.iter_start_state = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state11;
    assign seq_loop_intf_41.iter_end_state0 = AESL_inst_keygen.grp_iFFT_fu_1345.ap_ST_fsm_state13;
    assign seq_loop_intf_41.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_41.iter_end_state1 = 13'h0;
    assign seq_loop_intf_41.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_41.one_state_loop = 1'b0;
    assign seq_loop_intf_41.one_state_block = 1'b0;
    assign seq_loop_intf_41.finish = finish;
    csv_file_dump seq_loop_csv_dumper_41;
    seq_loop_monitor #(13) seq_loop_monitor_41;
    seq_loop_intf#(116) seq_loop_intf_42(clock,reset);
    assign seq_loop_intf_42.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state1;
    assign seq_loop_intf_42.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_42.pre_loop_state1 = 116'h0;
    assign seq_loop_intf_42.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_42.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state4;
    assign seq_loop_intf_42.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_42.post_loop_state1 = 116'h0;
    assign seq_loop_intf_42.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_42.post_loop_state2 = 116'h0;
    assign seq_loop_intf_42.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_42.post_loop_state3 = 116'h0;
    assign seq_loop_intf_42.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_42.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state2;
    assign seq_loop_intf_42.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_42.quit_loop_state1 = 116'h0;
    assign seq_loop_intf_42.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_42.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_CS_fsm;
    assign seq_loop_intf_42.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state2;
    assign seq_loop_intf_42.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state3;
    assign seq_loop_intf_42.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_42.iter_end_state1 = 116'h0;
    assign seq_loop_intf_42.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_42.one_state_loop = 1'b0;
    assign seq_loop_intf_42.one_state_block = 1'b0;
    assign seq_loop_intf_42.finish = finish;
    csv_file_dump seq_loop_csv_dumper_42;
    seq_loop_monitor #(116) seq_loop_monitor_42;
    seq_loop_intf#(116) seq_loop_intf_43(clock,reset);
    assign seq_loop_intf_43.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state4;
    assign seq_loop_intf_43.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_43.pre_loop_state1 = 116'h0;
    assign seq_loop_intf_43.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_43.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state97;
    assign seq_loop_intf_43.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_43.post_loop_state1 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state116;
    assign seq_loop_intf_43.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_43.post_loop_state2 = 116'h0;
    assign seq_loop_intf_43.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_43.post_loop_state3 = 116'h0;
    assign seq_loop_intf_43.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_43.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state5;
    assign seq_loop_intf_43.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_43.quit_loop_state1 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state6;
    assign seq_loop_intf_43.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_43.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_CS_fsm;
    assign seq_loop_intf_43.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state5;
    assign seq_loop_intf_43.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state96;
    assign seq_loop_intf_43.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_43.iter_end_state1 = 116'h0;
    assign seq_loop_intf_43.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_43.one_state_loop = 1'b0;
    assign seq_loop_intf_43.one_state_block = 1'b0;
    assign seq_loop_intf_43.finish = finish;
    csv_file_dump seq_loop_csv_dumper_43;
    seq_loop_monitor #(116) seq_loop_monitor_43;
    seq_loop_intf#(116) seq_loop_intf_44(clock,reset);
    assign seq_loop_intf_44.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state99;
    assign seq_loop_intf_44.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_44.pre_loop_state1 = 116'h0;
    assign seq_loop_intf_44.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_44.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state98;
    assign seq_loop_intf_44.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_44.post_loop_state1 = 116'h0;
    assign seq_loop_intf_44.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_44.post_loop_state2 = 116'h0;
    assign seq_loop_intf_44.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_44.post_loop_state3 = 116'h0;
    assign seq_loop_intf_44.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_44.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state100;
    assign seq_loop_intf_44.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_44.quit_loop_state1 = 116'h0;
    assign seq_loop_intf_44.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_44.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_CS_fsm;
    assign seq_loop_intf_44.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state100;
    assign seq_loop_intf_44.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state110;
    assign seq_loop_intf_44.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_44.iter_end_state1 = 116'h0;
    assign seq_loop_intf_44.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_44.one_state_loop = 1'b0;
    assign seq_loop_intf_44.one_state_block = 1'b0;
    assign seq_loop_intf_44.finish = finish;
    csv_file_dump seq_loop_csv_dumper_44;
    seq_loop_monitor #(116) seq_loop_monitor_44;
    seq_loop_intf#(116) seq_loop_intf_45(clock,reset);
    assign seq_loop_intf_45.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state97;
    assign seq_loop_intf_45.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_45.pre_loop_state1 = 116'h0;
    assign seq_loop_intf_45.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_45.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state97;
    assign seq_loop_intf_45.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_45.post_loop_state1 = 116'h0;
    assign seq_loop_intf_45.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_45.post_loop_state2 = 116'h0;
    assign seq_loop_intf_45.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_45.post_loop_state3 = 116'h0;
    assign seq_loop_intf_45.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_45.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state98;
    assign seq_loop_intf_45.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_45.quit_loop_state1 = 116'h0;
    assign seq_loop_intf_45.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_45.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_CS_fsm;
    assign seq_loop_intf_45.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state98;
    assign seq_loop_intf_45.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state100;
    assign seq_loop_intf_45.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_45.iter_end_state1 = 116'h0;
    assign seq_loop_intf_45.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_45.one_state_loop = 1'b0;
    assign seq_loop_intf_45.one_state_block = 1'b0;
    assign seq_loop_intf_45.finish = finish;
    csv_file_dump seq_loop_csv_dumper_45;
    seq_loop_monitor #(116) seq_loop_monitor_45;
    seq_loop_intf#(116) seq_loop_intf_46(clock,reset);
    assign seq_loop_intf_46.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state5;
    assign seq_loop_intf_46.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_46.pre_loop_state1 = 116'h0;
    assign seq_loop_intf_46.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_46.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state111;
    assign seq_loop_intf_46.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_46.post_loop_state1 = 116'h0;
    assign seq_loop_intf_46.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_46.post_loop_state2 = 116'h0;
    assign seq_loop_intf_46.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_46.post_loop_state3 = 116'h0;
    assign seq_loop_intf_46.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_46.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state97;
    assign seq_loop_intf_46.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_46.quit_loop_state1 = 116'h0;
    assign seq_loop_intf_46.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_46.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_CS_fsm;
    assign seq_loop_intf_46.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state97;
    assign seq_loop_intf_46.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state98;
    assign seq_loop_intf_46.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_46.iter_end_state1 = 116'h0;
    assign seq_loop_intf_46.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_46.one_state_loop = 1'b0;
    assign seq_loop_intf_46.one_state_block = 1'b0;
    assign seq_loop_intf_46.finish = finish;
    csv_file_dump seq_loop_csv_dumper_46;
    seq_loop_monitor #(116) seq_loop_monitor_46;
    seq_loop_intf#(116) seq_loop_intf_47(clock,reset);
    assign seq_loop_intf_47.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state97;
    assign seq_loop_intf_47.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_47.pre_loop_state1 = 116'h0;
    assign seq_loop_intf_47.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_47.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state116;
    assign seq_loop_intf_47.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_47.post_loop_state1 = 116'h0;
    assign seq_loop_intf_47.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_47.post_loop_state2 = 116'h0;
    assign seq_loop_intf_47.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_47.post_loop_state3 = 116'h0;
    assign seq_loop_intf_47.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_47.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state111;
    assign seq_loop_intf_47.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_47.quit_loop_state1 = 116'h0;
    assign seq_loop_intf_47.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_47.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_CS_fsm;
    assign seq_loop_intf_47.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state111;
    assign seq_loop_intf_47.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.ap_ST_fsm_state115;
    assign seq_loop_intf_47.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_47.iter_end_state1 = 116'h0;
    assign seq_loop_intf_47.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_47.one_state_loop = 1'b0;
    assign seq_loop_intf_47.one_state_block = 1'b0;
    assign seq_loop_intf_47.finish = finish;
    csv_file_dump seq_loop_csv_dumper_47;
    seq_loop_monitor #(116) seq_loop_monitor_47;
    seq_loop_intf#(16) seq_loop_intf_48(clock,reset);
    assign seq_loop_intf_48.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state4;
    assign seq_loop_intf_48.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_48.pre_loop_state1 = 16'h0;
    assign seq_loop_intf_48.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_48.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state3;
    assign seq_loop_intf_48.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_48.post_loop_state1 = 16'h0;
    assign seq_loop_intf_48.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_48.post_loop_state2 = 16'h0;
    assign seq_loop_intf_48.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_48.post_loop_state3 = 16'h0;
    assign seq_loop_intf_48.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_48.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state5;
    assign seq_loop_intf_48.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_48.quit_loop_state1 = 16'h0;
    assign seq_loop_intf_48.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_48.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_CS_fsm;
    assign seq_loop_intf_48.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state5;
    assign seq_loop_intf_48.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state16;
    assign seq_loop_intf_48.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_48.iter_end_state1 = 16'h0;
    assign seq_loop_intf_48.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_48.one_state_loop = 1'b0;
    assign seq_loop_intf_48.one_state_block = 1'b0;
    assign seq_loop_intf_48.finish = finish;
    csv_file_dump seq_loop_csv_dumper_48;
    seq_loop_monitor #(16) seq_loop_monitor_48;
    seq_loop_intf#(16) seq_loop_intf_49(clock,reset);
    assign seq_loop_intf_49.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state2;
    assign seq_loop_intf_49.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_49.pre_loop_state1 = 16'h0;
    assign seq_loop_intf_49.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_49.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state2;
    assign seq_loop_intf_49.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_49.post_loop_state1 = 16'h0;
    assign seq_loop_intf_49.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_49.post_loop_state2 = 16'h0;
    assign seq_loop_intf_49.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_49.post_loop_state3 = 16'h0;
    assign seq_loop_intf_49.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_49.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state3;
    assign seq_loop_intf_49.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_49.quit_loop_state1 = 16'h0;
    assign seq_loop_intf_49.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_49.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_CS_fsm;
    assign seq_loop_intf_49.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state3;
    assign seq_loop_intf_49.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state5;
    assign seq_loop_intf_49.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_49.iter_end_state1 = 16'h0;
    assign seq_loop_intf_49.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_49.one_state_loop = 1'b0;
    assign seq_loop_intf_49.one_state_block = 1'b0;
    assign seq_loop_intf_49.finish = finish;
    csv_file_dump seq_loop_csv_dumper_49;
    seq_loop_monitor #(16) seq_loop_monitor_49;
    seq_loop_intf#(16) seq_loop_intf_50(clock,reset);
    assign seq_loop_intf_50.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state1;
    assign seq_loop_intf_50.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_50.pre_loop_state1 = 16'h0;
    assign seq_loop_intf_50.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_50.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state1;
    assign seq_loop_intf_50.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_50.post_loop_state1 = 16'h0;
    assign seq_loop_intf_50.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_50.post_loop_state2 = 16'h0;
    assign seq_loop_intf_50.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_50.post_loop_state3 = 16'h0;
    assign seq_loop_intf_50.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_50.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state2;
    assign seq_loop_intf_50.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_50.quit_loop_state1 = 16'h0;
    assign seq_loop_intf_50.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_50.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_CS_fsm;
    assign seq_loop_intf_50.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state2;
    assign seq_loop_intf_50.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_fu_320.ap_ST_fsm_state3;
    assign seq_loop_intf_50.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_50.iter_end_state1 = 16'h0;
    assign seq_loop_intf_50.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_50.one_state_loop = 1'b0;
    assign seq_loop_intf_50.one_state_block = 1'b0;
    assign seq_loop_intf_50.finish = finish;
    csv_file_dump seq_loop_csv_dumper_50;
    seq_loop_monitor #(16) seq_loop_monitor_50;
    seq_loop_intf#(16) seq_loop_intf_51(clock,reset);
    assign seq_loop_intf_51.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state4;
    assign seq_loop_intf_51.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_51.pre_loop_state1 = 16'h0;
    assign seq_loop_intf_51.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_51.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state3;
    assign seq_loop_intf_51.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_51.post_loop_state1 = 16'h0;
    assign seq_loop_intf_51.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_51.post_loop_state2 = 16'h0;
    assign seq_loop_intf_51.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_51.post_loop_state3 = 16'h0;
    assign seq_loop_intf_51.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_51.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state5;
    assign seq_loop_intf_51.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_51.quit_loop_state1 = 16'h0;
    assign seq_loop_intf_51.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_51.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_CS_fsm;
    assign seq_loop_intf_51.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state5;
    assign seq_loop_intf_51.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state16;
    assign seq_loop_intf_51.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_51.iter_end_state1 = 16'h0;
    assign seq_loop_intf_51.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_51.one_state_loop = 1'b0;
    assign seq_loop_intf_51.one_state_block = 1'b0;
    assign seq_loop_intf_51.finish = finish;
    csv_file_dump seq_loop_csv_dumper_51;
    seq_loop_monitor #(16) seq_loop_monitor_51;
    seq_loop_intf#(16) seq_loop_intf_52(clock,reset);
    assign seq_loop_intf_52.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state2;
    assign seq_loop_intf_52.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_52.pre_loop_state1 = 16'h0;
    assign seq_loop_intf_52.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_52.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state2;
    assign seq_loop_intf_52.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_52.post_loop_state1 = 16'h0;
    assign seq_loop_intf_52.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_52.post_loop_state2 = 16'h0;
    assign seq_loop_intf_52.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_52.post_loop_state3 = 16'h0;
    assign seq_loop_intf_52.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_52.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state3;
    assign seq_loop_intf_52.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_52.quit_loop_state1 = 16'h0;
    assign seq_loop_intf_52.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_52.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_CS_fsm;
    assign seq_loop_intf_52.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state3;
    assign seq_loop_intf_52.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state5;
    assign seq_loop_intf_52.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_52.iter_end_state1 = 16'h0;
    assign seq_loop_intf_52.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_52.one_state_loop = 1'b0;
    assign seq_loop_intf_52.one_state_block = 1'b0;
    assign seq_loop_intf_52.finish = finish;
    csv_file_dump seq_loop_csv_dumper_52;
    seq_loop_monitor #(16) seq_loop_monitor_52;
    seq_loop_intf#(16) seq_loop_intf_53(clock,reset);
    assign seq_loop_intf_53.pre_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state1;
    assign seq_loop_intf_53.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_53.pre_loop_state1 = 16'h0;
    assign seq_loop_intf_53.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_53.post_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state1;
    assign seq_loop_intf_53.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_53.post_loop_state1 = 16'h0;
    assign seq_loop_intf_53.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_53.post_loop_state2 = 16'h0;
    assign seq_loop_intf_53.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_53.post_loop_state3 = 16'h0;
    assign seq_loop_intf_53.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_53.quit_loop_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state2;
    assign seq_loop_intf_53.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_53.quit_loop_state1 = 16'h0;
    assign seq_loop_intf_53.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_53.cur_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_CS_fsm;
    assign seq_loop_intf_53.iter_start_state = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state2;
    assign seq_loop_intf_53.iter_end_state0 = AESL_inst_keygen.grp_compute_public_1_fu_1352.grp_mq_NTT_1_fu_328.ap_ST_fsm_state3;
    assign seq_loop_intf_53.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_53.iter_end_state1 = 16'h0;
    assign seq_loop_intf_53.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_53.one_state_loop = 1'b0;
    assign seq_loop_intf_53.one_state_block = 1'b0;
    assign seq_loop_intf_53.finish = finish;
    csv_file_dump seq_loop_csv_dumper_53;
    seq_loop_monitor #(16) seq_loop_monitor_53;
    seq_loop_intf#(31) seq_loop_intf_54(clock,reset);
    assign seq_loop_intf_54.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state2;
    assign seq_loop_intf_54.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_54.pre_loop_state1 = 31'h0;
    assign seq_loop_intf_54.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_54.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state5;
    assign seq_loop_intf_54.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_54.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state31;
    assign seq_loop_intf_54.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_54.post_loop_state2 = 31'h0;
    assign seq_loop_intf_54.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_54.post_loop_state3 = 31'h0;
    assign seq_loop_intf_54.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_54.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state4;
    assign seq_loop_intf_54.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_54.quit_loop_state1 = 31'h0;
    assign seq_loop_intf_54.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_54.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_CS_fsm;
    assign seq_loop_intf_54.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state3;
    assign seq_loop_intf_54.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state4;
    assign seq_loop_intf_54.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_54.iter_end_state1 = 31'h0;
    assign seq_loop_intf_54.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_54.one_state_loop = 1'b0;
    assign seq_loop_intf_54.one_state_block = 1'b0;
    assign seq_loop_intf_54.finish = finish;
    csv_file_dump seq_loop_csv_dumper_54;
    seq_loop_monitor #(31) seq_loop_monitor_54;
    seq_loop_intf#(31) seq_loop_intf_55(clock,reset);
    assign seq_loop_intf_55.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state8;
    assign seq_loop_intf_55.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_55.pre_loop_state1 = 31'h0;
    assign seq_loop_intf_55.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_55.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state11;
    assign seq_loop_intf_55.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_55.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state12;
    assign seq_loop_intf_55.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_55.post_loop_state2 = 31'h0;
    assign seq_loop_intf_55.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_55.post_loop_state3 = 31'h0;
    assign seq_loop_intf_55.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_55.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state9;
    assign seq_loop_intf_55.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_55.quit_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state10;
    assign seq_loop_intf_55.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_55.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_CS_fsm;
    assign seq_loop_intf_55.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state9;
    assign seq_loop_intf_55.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state10;
    assign seq_loop_intf_55.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_55.iter_end_state1 = 31'h0;
    assign seq_loop_intf_55.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_55.one_state_loop = 1'b0;
    assign seq_loop_intf_55.one_state_block = 1'b0;
    assign seq_loop_intf_55.finish = finish;
    csv_file_dump seq_loop_csv_dumper_55;
    seq_loop_monitor #(31) seq_loop_monitor_55;
    seq_loop_intf#(31) seq_loop_intf_56(clock,reset);
    assign seq_loop_intf_56.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state9;
    assign seq_loop_intf_56.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_56.pre_loop_state1 = 31'h0;
    assign seq_loop_intf_56.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_56.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state13;
    assign seq_loop_intf_56.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_56.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state31;
    assign seq_loop_intf_56.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_56.post_loop_state2 = 31'h0;
    assign seq_loop_intf_56.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_56.post_loop_state3 = 31'h0;
    assign seq_loop_intf_56.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_56.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state11;
    assign seq_loop_intf_56.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_56.quit_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state12;
    assign seq_loop_intf_56.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_56.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_CS_fsm;
    assign seq_loop_intf_56.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state11;
    assign seq_loop_intf_56.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state12;
    assign seq_loop_intf_56.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_56.iter_end_state1 = 31'h0;
    assign seq_loop_intf_56.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_56.one_state_loop = 1'b0;
    assign seq_loop_intf_56.one_state_block = 1'b0;
    assign seq_loop_intf_56.finish = finish;
    csv_file_dump seq_loop_csv_dumper_56;
    seq_loop_monitor #(31) seq_loop_monitor_56;
    seq_loop_intf#(31) seq_loop_intf_57(clock,reset);
    assign seq_loop_intf_57.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state11;
    assign seq_loop_intf_57.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_57.pre_loop_state1 = 31'h0;
    assign seq_loop_intf_57.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_57.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state15;
    assign seq_loop_intf_57.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_57.post_loop_state1 = 31'h0;
    assign seq_loop_intf_57.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_57.post_loop_state2 = 31'h0;
    assign seq_loop_intf_57.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_57.post_loop_state3 = 31'h0;
    assign seq_loop_intf_57.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_57.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state13;
    assign seq_loop_intf_57.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_57.quit_loop_state1 = 31'h0;
    assign seq_loop_intf_57.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_57.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_CS_fsm;
    assign seq_loop_intf_57.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state13;
    assign seq_loop_intf_57.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state14;
    assign seq_loop_intf_57.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_57.iter_end_state1 = 31'h0;
    assign seq_loop_intf_57.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_57.one_state_loop = 1'b0;
    assign seq_loop_intf_57.one_state_block = 1'b0;
    assign seq_loop_intf_57.finish = finish;
    csv_file_dump seq_loop_csv_dumper_57;
    seq_loop_monitor #(31) seq_loop_monitor_57;
    seq_loop_intf#(31) seq_loop_intf_58(clock,reset);
    assign seq_loop_intf_58.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state13;
    assign seq_loop_intf_58.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_58.pre_loop_state1 = 31'h0;
    assign seq_loop_intf_58.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_58.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state17;
    assign seq_loop_intf_58.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_58.post_loop_state1 = 31'h0;
    assign seq_loop_intf_58.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_58.post_loop_state2 = 31'h0;
    assign seq_loop_intf_58.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_58.post_loop_state3 = 31'h0;
    assign seq_loop_intf_58.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_58.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state15;
    assign seq_loop_intf_58.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_58.quit_loop_state1 = 31'h0;
    assign seq_loop_intf_58.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_58.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_CS_fsm;
    assign seq_loop_intf_58.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state15;
    assign seq_loop_intf_58.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state16;
    assign seq_loop_intf_58.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_58.iter_end_state1 = 31'h0;
    assign seq_loop_intf_58.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_58.one_state_loop = 1'b0;
    assign seq_loop_intf_58.one_state_block = 1'b0;
    assign seq_loop_intf_58.finish = finish;
    csv_file_dump seq_loop_csv_dumper_58;
    seq_loop_monitor #(31) seq_loop_monitor_58;
    seq_loop_intf#(31) seq_loop_intf_59(clock,reset);
    assign seq_loop_intf_59.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state15;
    assign seq_loop_intf_59.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_59.pre_loop_state1 = 31'h0;
    assign seq_loop_intf_59.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_59.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state19;
    assign seq_loop_intf_59.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_59.post_loop_state1 = 31'h0;
    assign seq_loop_intf_59.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_59.post_loop_state2 = 31'h0;
    assign seq_loop_intf_59.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_59.post_loop_state3 = 31'h0;
    assign seq_loop_intf_59.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_59.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state17;
    assign seq_loop_intf_59.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_59.quit_loop_state1 = 31'h0;
    assign seq_loop_intf_59.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_59.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_CS_fsm;
    assign seq_loop_intf_59.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state17;
    assign seq_loop_intf_59.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state18;
    assign seq_loop_intf_59.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_59.iter_end_state1 = 31'h0;
    assign seq_loop_intf_59.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_59.one_state_loop = 1'b0;
    assign seq_loop_intf_59.one_state_block = 1'b0;
    assign seq_loop_intf_59.finish = finish;
    csv_file_dump seq_loop_csv_dumper_59;
    seq_loop_monitor #(31) seq_loop_monitor_59;
    seq_loop_intf#(31) seq_loop_intf_60(clock,reset);
    assign seq_loop_intf_60.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state17;
    assign seq_loop_intf_60.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_60.pre_loop_state1 = 31'h0;
    assign seq_loop_intf_60.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_60.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state22;
    assign seq_loop_intf_60.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_60.post_loop_state1 = 31'h0;
    assign seq_loop_intf_60.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_60.post_loop_state2 = 31'h0;
    assign seq_loop_intf_60.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_60.post_loop_state3 = 31'h0;
    assign seq_loop_intf_60.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_60.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state19;
    assign seq_loop_intf_60.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_60.quit_loop_state1 = 31'h0;
    assign seq_loop_intf_60.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_60.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_CS_fsm;
    assign seq_loop_intf_60.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state19;
    assign seq_loop_intf_60.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state21;
    assign seq_loop_intf_60.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_60.iter_end_state1 = 31'h0;
    assign seq_loop_intf_60.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_60.one_state_loop = 1'b0;
    assign seq_loop_intf_60.one_state_block = 1'b0;
    assign seq_loop_intf_60.finish = finish;
    csv_file_dump seq_loop_csv_dumper_60;
    seq_loop_monitor #(31) seq_loop_monitor_60;
    seq_loop_intf#(31) seq_loop_intf_61(clock,reset);
    assign seq_loop_intf_61.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state28;
    assign seq_loop_intf_61.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_61.pre_loop_state1 = 31'h0;
    assign seq_loop_intf_61.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_61.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state1;
    assign seq_loop_intf_61.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_61.post_loop_state1 = 31'h0;
    assign seq_loop_intf_61.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_61.post_loop_state2 = 31'h0;
    assign seq_loop_intf_61.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_61.post_loop_state3 = 31'h0;
    assign seq_loop_intf_61.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_61.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state29;
    assign seq_loop_intf_61.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_61.quit_loop_state1 = 31'h0;
    assign seq_loop_intf_61.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_61.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_CS_fsm;
    assign seq_loop_intf_61.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state29;
    assign seq_loop_intf_61.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.ap_ST_fsm_state31;
    assign seq_loop_intf_61.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_61.iter_end_state1 = 31'h0;
    assign seq_loop_intf_61.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_61.one_state_loop = 1'b0;
    assign seq_loop_intf_61.one_state_block = 1'b0;
    assign seq_loop_intf_61.finish = finish;
    csv_file_dump seq_loop_csv_dumper_61;
    seq_loop_monitor #(31) seq_loop_monitor_61;
    seq_loop_intf#(452) seq_loop_intf_62(clock,reset);
    assign seq_loop_intf_62.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state269;
    assign seq_loop_intf_62.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_62.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_62.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_62.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state272;
    assign seq_loop_intf_62.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_62.post_loop_state1 = 452'h0;
    assign seq_loop_intf_62.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_62.post_loop_state2 = 452'h0;
    assign seq_loop_intf_62.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_62.post_loop_state3 = 452'h0;
    assign seq_loop_intf_62.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_62.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state270;
    assign seq_loop_intf_62.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_62.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_62.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_62.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_62.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state270;
    assign seq_loop_intf_62.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state271;
    assign seq_loop_intf_62.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_62.iter_end_state1 = 452'h0;
    assign seq_loop_intf_62.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_62.one_state_loop = 1'b0;
    assign seq_loop_intf_62.one_state_block = 1'b0;
    assign seq_loop_intf_62.finish = finish;
    csv_file_dump seq_loop_csv_dumper_62;
    seq_loop_monitor #(452) seq_loop_monitor_62;
    seq_loop_intf#(452) seq_loop_intf_63(clock,reset);
    assign seq_loop_intf_63.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state270;
    assign seq_loop_intf_63.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_63.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_63.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_63.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state452;
    assign seq_loop_intf_63.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_63.post_loop_state1 = 452'h0;
    assign seq_loop_intf_63.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_63.post_loop_state2 = 452'h0;
    assign seq_loop_intf_63.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_63.post_loop_state3 = 452'h0;
    assign seq_loop_intf_63.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_63.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state272;
    assign seq_loop_intf_63.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_63.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_63.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_63.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_63.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state272;
    assign seq_loop_intf_63.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state273;
    assign seq_loop_intf_63.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_63.iter_end_state1 = 452'h0;
    assign seq_loop_intf_63.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_63.one_state_loop = 1'b0;
    assign seq_loop_intf_63.one_state_block = 1'b0;
    assign seq_loop_intf_63.finish = finish;
    csv_file_dump seq_loop_csv_dumper_63;
    seq_loop_monitor #(452) seq_loop_monitor_63;
    seq_loop_intf#(452) seq_loop_intf_64(clock,reset);
    assign seq_loop_intf_64.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state110;
    assign seq_loop_intf_64.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_64.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_64.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_64.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state113;
    assign seq_loop_intf_64.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_64.post_loop_state1 = 452'h0;
    assign seq_loop_intf_64.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_64.post_loop_state2 = 452'h0;
    assign seq_loop_intf_64.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_64.post_loop_state3 = 452'h0;
    assign seq_loop_intf_64.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_64.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state111;
    assign seq_loop_intf_64.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_64.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_64.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_64.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_64.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state111;
    assign seq_loop_intf_64.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state112;
    assign seq_loop_intf_64.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_64.iter_end_state1 = 452'h0;
    assign seq_loop_intf_64.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_64.one_state_loop = 1'b0;
    assign seq_loop_intf_64.one_state_block = 1'b0;
    assign seq_loop_intf_64.finish = finish;
    csv_file_dump seq_loop_csv_dumper_64;
    seq_loop_monitor #(452) seq_loop_monitor_64;
    seq_loop_intf#(452) seq_loop_intf_65(clock,reset);
    assign seq_loop_intf_65.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state111;
    assign seq_loop_intf_65.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_65.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_65.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_65.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state106;
    assign seq_loop_intf_65.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_65.post_loop_state1 = 452'h0;
    assign seq_loop_intf_65.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_65.post_loop_state2 = 452'h0;
    assign seq_loop_intf_65.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_65.post_loop_state3 = 452'h0;
    assign seq_loop_intf_65.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_65.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state113;
    assign seq_loop_intf_65.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_65.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_65.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_65.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_65.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state113;
    assign seq_loop_intf_65.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state118;
    assign seq_loop_intf_65.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_65.iter_end_state1 = 452'h0;
    assign seq_loop_intf_65.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_65.one_state_loop = 1'b0;
    assign seq_loop_intf_65.one_state_block = 1'b0;
    assign seq_loop_intf_65.finish = finish;
    csv_file_dump seq_loop_csv_dumper_65;
    seq_loop_monitor #(452) seq_loop_monitor_65;
    seq_loop_intf#(452) seq_loop_intf_66(clock,reset);
    assign seq_loop_intf_66.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state1;
    assign seq_loop_intf_66.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_66.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_66.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_66.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state119;
    assign seq_loop_intf_66.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_66.post_loop_state1 = 452'h0;
    assign seq_loop_intf_66.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_66.post_loop_state2 = 452'h0;
    assign seq_loop_intf_66.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_66.post_loop_state3 = 452'h0;
    assign seq_loop_intf_66.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_66.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state106;
    assign seq_loop_intf_66.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_66.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_66.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_66.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_66.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state106;
    assign seq_loop_intf_66.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state113;
    assign seq_loop_intf_66.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_66.iter_end_state1 = 452'h0;
    assign seq_loop_intf_66.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_66.one_state_loop = 1'b0;
    assign seq_loop_intf_66.one_state_block = 1'b0;
    assign seq_loop_intf_66.finish = finish;
    csv_file_dump seq_loop_csv_dumper_66;
    seq_loop_monitor #(452) seq_loop_monitor_66;
    seq_loop_intf#(452) seq_loop_intf_67(clock,reset);
    assign seq_loop_intf_67.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state106;
    assign seq_loop_intf_67.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_67.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_67.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_67.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state121;
    assign seq_loop_intf_67.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_67.post_loop_state1 = 452'h0;
    assign seq_loop_intf_67.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_67.post_loop_state2 = 452'h0;
    assign seq_loop_intf_67.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_67.post_loop_state3 = 452'h0;
    assign seq_loop_intf_67.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_67.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state120;
    assign seq_loop_intf_67.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_67.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_67.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_67.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_67.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state119;
    assign seq_loop_intf_67.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state120;
    assign seq_loop_intf_67.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_67.iter_end_state1 = 452'h0;
    assign seq_loop_intf_67.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_67.one_state_loop = 1'b0;
    assign seq_loop_intf_67.one_state_block = 1'b0;
    assign seq_loop_intf_67.finish = finish;
    csv_file_dump seq_loop_csv_dumper_67;
    seq_loop_monitor #(452) seq_loop_monitor_67;
    seq_loop_intf#(452) seq_loop_intf_68(clock,reset);
    assign seq_loop_intf_68.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state120;
    assign seq_loop_intf_68.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_68.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_68.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_68.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state123;
    assign seq_loop_intf_68.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_68.post_loop_state1 = 452'h0;
    assign seq_loop_intf_68.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_68.post_loop_state2 = 452'h0;
    assign seq_loop_intf_68.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_68.post_loop_state3 = 452'h0;
    assign seq_loop_intf_68.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_68.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state122;
    assign seq_loop_intf_68.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_68.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_68.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_68.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_68.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state121;
    assign seq_loop_intf_68.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state122;
    assign seq_loop_intf_68.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_68.iter_end_state1 = 452'h0;
    assign seq_loop_intf_68.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_68.one_state_loop = 1'b0;
    assign seq_loop_intf_68.one_state_block = 1'b0;
    assign seq_loop_intf_68.finish = finish;
    csv_file_dump seq_loop_csv_dumper_68;
    seq_loop_monitor #(452) seq_loop_monitor_68;
    seq_loop_intf#(452) seq_loop_intf_69(clock,reset);
    assign seq_loop_intf_69.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state127;
    assign seq_loop_intf_69.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_69.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_69.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_69.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state130;
    assign seq_loop_intf_69.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_69.post_loop_state1 = 452'h0;
    assign seq_loop_intf_69.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_69.post_loop_state2 = 452'h0;
    assign seq_loop_intf_69.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_69.post_loop_state3 = 452'h0;
    assign seq_loop_intf_69.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_69.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state128;
    assign seq_loop_intf_69.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_69.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_69.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_69.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_69.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state128;
    assign seq_loop_intf_69.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state129;
    assign seq_loop_intf_69.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_69.iter_end_state1 = 452'h0;
    assign seq_loop_intf_69.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_69.one_state_loop = 1'b0;
    assign seq_loop_intf_69.one_state_block = 1'b0;
    assign seq_loop_intf_69.finish = finish;
    csv_file_dump seq_loop_csv_dumper_69;
    seq_loop_monitor #(452) seq_loop_monitor_69;
    seq_loop_intf#(452) seq_loop_intf_70(clock,reset);
    assign seq_loop_intf_70.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state132;
    assign seq_loop_intf_70.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_70.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_70.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_70.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state136;
    assign seq_loop_intf_70.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_70.post_loop_state1 = 452'h0;
    assign seq_loop_intf_70.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_70.post_loop_state2 = 452'h0;
    assign seq_loop_intf_70.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_70.post_loop_state3 = 452'h0;
    assign seq_loop_intf_70.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_70.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state133;
    assign seq_loop_intf_70.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_70.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_70.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_70.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_70.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state133;
    assign seq_loop_intf_70.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state135;
    assign seq_loop_intf_70.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_70.iter_end_state1 = 452'h0;
    assign seq_loop_intf_70.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_70.one_state_loop = 1'b0;
    assign seq_loop_intf_70.one_state_block = 1'b0;
    assign seq_loop_intf_70.finish = finish;
    csv_file_dump seq_loop_csv_dumper_70;
    seq_loop_monitor #(452) seq_loop_monitor_70;
    seq_loop_intf#(452) seq_loop_intf_71(clock,reset);
    assign seq_loop_intf_71.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state133;
    assign seq_loop_intf_71.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_71.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_71.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_71.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state139;
    assign seq_loop_intf_71.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_71.post_loop_state1 = 452'h0;
    assign seq_loop_intf_71.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_71.post_loop_state2 = 452'h0;
    assign seq_loop_intf_71.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_71.post_loop_state3 = 452'h0;
    assign seq_loop_intf_71.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_71.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state136;
    assign seq_loop_intf_71.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_71.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_71.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_71.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_71.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state136;
    assign seq_loop_intf_71.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state138;
    assign seq_loop_intf_71.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_71.iter_end_state1 = 452'h0;
    assign seq_loop_intf_71.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_71.one_state_loop = 1'b0;
    assign seq_loop_intf_71.one_state_block = 1'b0;
    assign seq_loop_intf_71.finish = finish;
    csv_file_dump seq_loop_csv_dumper_71;
    seq_loop_monitor #(452) seq_loop_monitor_71;
    seq_loop_intf#(452) seq_loop_intf_72(clock,reset);
    assign seq_loop_intf_72.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state136;
    assign seq_loop_intf_72.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_72.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_72.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_72.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state141;
    assign seq_loop_intf_72.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_72.post_loop_state1 = 452'h0;
    assign seq_loop_intf_72.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_72.post_loop_state2 = 452'h0;
    assign seq_loop_intf_72.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_72.post_loop_state3 = 452'h0;
    assign seq_loop_intf_72.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_72.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state140;
    assign seq_loop_intf_72.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_72.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_72.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_72.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_72.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state139;
    assign seq_loop_intf_72.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state140;
    assign seq_loop_intf_72.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_72.iter_end_state1 = 452'h0;
    assign seq_loop_intf_72.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_72.one_state_loop = 1'b0;
    assign seq_loop_intf_72.one_state_block = 1'b0;
    assign seq_loop_intf_72.finish = finish;
    csv_file_dump seq_loop_csv_dumper_72;
    seq_loop_monitor #(452) seq_loop_monitor_72;
    seq_loop_intf#(452) seq_loop_intf_73(clock,reset);
    assign seq_loop_intf_73.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state140;
    assign seq_loop_intf_73.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_73.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_73.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_73.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state143;
    assign seq_loop_intf_73.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_73.post_loop_state1 = 452'h0;
    assign seq_loop_intf_73.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_73.post_loop_state2 = 452'h0;
    assign seq_loop_intf_73.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_73.post_loop_state3 = 452'h0;
    assign seq_loop_intf_73.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_73.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state142;
    assign seq_loop_intf_73.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_73.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_73.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_73.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_73.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state141;
    assign seq_loop_intf_73.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state142;
    assign seq_loop_intf_73.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_73.iter_end_state1 = 452'h0;
    assign seq_loop_intf_73.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_73.one_state_loop = 1'b0;
    assign seq_loop_intf_73.one_state_block = 1'b0;
    assign seq_loop_intf_73.finish = finish;
    csv_file_dump seq_loop_csv_dumper_73;
    seq_loop_monitor #(452) seq_loop_monitor_73;
    seq_loop_intf#(452) seq_loop_intf_74(clock,reset);
    assign seq_loop_intf_74.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state142;
    assign seq_loop_intf_74.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_74.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_74.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_74.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state145;
    assign seq_loop_intf_74.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_74.post_loop_state1 = 452'h0;
    assign seq_loop_intf_74.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_74.post_loop_state2 = 452'h0;
    assign seq_loop_intf_74.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_74.post_loop_state3 = 452'h0;
    assign seq_loop_intf_74.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_74.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state144;
    assign seq_loop_intf_74.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_74.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_74.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_74.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_74.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state143;
    assign seq_loop_intf_74.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state144;
    assign seq_loop_intf_74.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_74.iter_end_state1 = 452'h0;
    assign seq_loop_intf_74.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_74.one_state_loop = 1'b0;
    assign seq_loop_intf_74.one_state_block = 1'b0;
    assign seq_loop_intf_74.finish = finish;
    csv_file_dump seq_loop_csv_dumper_74;
    seq_loop_monitor #(452) seq_loop_monitor_74;
    seq_loop_intf#(452) seq_loop_intf_75(clock,reset);
    assign seq_loop_intf_75.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state144;
    assign seq_loop_intf_75.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_75.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_75.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_75.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state149;
    assign seq_loop_intf_75.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_75.post_loop_state1 = 452'h0;
    assign seq_loop_intf_75.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_75.post_loop_state2 = 452'h0;
    assign seq_loop_intf_75.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_75.post_loop_state3 = 452'h0;
    assign seq_loop_intf_75.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_75.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state145;
    assign seq_loop_intf_75.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_75.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_75.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_75.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_75.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state145;
    assign seq_loop_intf_75.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state148;
    assign seq_loop_intf_75.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_75.iter_end_state1 = 452'h0;
    assign seq_loop_intf_75.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_75.one_state_loop = 1'b0;
    assign seq_loop_intf_75.one_state_block = 1'b0;
    assign seq_loop_intf_75.finish = finish;
    csv_file_dump seq_loop_csv_dumper_75;
    seq_loop_monitor #(452) seq_loop_monitor_75;
    seq_loop_intf#(452) seq_loop_intf_76(clock,reset);
    assign seq_loop_intf_76.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state151;
    assign seq_loop_intf_76.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_76.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_76.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_76.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state159;
    assign seq_loop_intf_76.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_76.post_loop_state1 = 452'h0;
    assign seq_loop_intf_76.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_76.post_loop_state2 = 452'h0;
    assign seq_loop_intf_76.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_76.post_loop_state3 = 452'h0;
    assign seq_loop_intf_76.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_76.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state152;
    assign seq_loop_intf_76.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_76.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_76.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_76.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_76.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state152;
    assign seq_loop_intf_76.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state158;
    assign seq_loop_intf_76.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_76.iter_end_state1 = 452'h0;
    assign seq_loop_intf_76.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_76.one_state_loop = 1'b0;
    assign seq_loop_intf_76.one_state_block = 1'b0;
    assign seq_loop_intf_76.finish = finish;
    csv_file_dump seq_loop_csv_dumper_76;
    seq_loop_monitor #(452) seq_loop_monitor_76;
    seq_loop_intf#(452) seq_loop_intf_77(clock,reset);
    assign seq_loop_intf_77.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state161;
    assign seq_loop_intf_77.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_77.pre_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state165;
    assign seq_loop_intf_77.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_77.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state123;
    assign seq_loop_intf_77.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_77.post_loop_state1 = 452'h0;
    assign seq_loop_intf_77.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_77.post_loop_state2 = 452'h0;
    assign seq_loop_intf_77.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_77.post_loop_state3 = 452'h0;
    assign seq_loop_intf_77.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_77.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state166;
    assign seq_loop_intf_77.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_77.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_77.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_77.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_77.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state166;
    assign seq_loop_intf_77.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state167;
    assign seq_loop_intf_77.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_77.iter_end_state1 = 452'h0;
    assign seq_loop_intf_77.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_77.one_state_loop = 1'b0;
    assign seq_loop_intf_77.one_state_block = 1'b0;
    assign seq_loop_intf_77.finish = finish;
    csv_file_dump seq_loop_csv_dumper_77;
    seq_loop_monitor #(452) seq_loop_monitor_77;
    seq_loop_intf#(452) seq_loop_intf_78(clock,reset);
    assign seq_loop_intf_78.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state122;
    assign seq_loop_intf_78.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_78.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_78.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_78.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state168;
    assign seq_loop_intf_78.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_78.post_loop_state1 = 452'h0;
    assign seq_loop_intf_78.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_78.post_loop_state2 = 452'h0;
    assign seq_loop_intf_78.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_78.post_loop_state3 = 452'h0;
    assign seq_loop_intf_78.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_78.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state123;
    assign seq_loop_intf_78.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_78.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_78.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_78.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_78.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state123;
    assign seq_loop_intf_78.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state166;
    assign seq_loop_intf_78.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_78.iter_end_state1 = 452'h0;
    assign seq_loop_intf_78.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_78.one_state_loop = 1'b0;
    assign seq_loop_intf_78.one_state_block = 1'b0;
    assign seq_loop_intf_78.finish = finish;
    csv_file_dump seq_loop_csv_dumper_78;
    seq_loop_monitor #(452) seq_loop_monitor_78;
    seq_loop_intf#(452) seq_loop_intf_79(clock,reset);
    assign seq_loop_intf_79.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state174;
    assign seq_loop_intf_79.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_79.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_79.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_79.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state177;
    assign seq_loop_intf_79.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_79.post_loop_state1 = 452'h0;
    assign seq_loop_intf_79.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_79.post_loop_state2 = 452'h0;
    assign seq_loop_intf_79.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_79.post_loop_state3 = 452'h0;
    assign seq_loop_intf_79.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_79.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state176;
    assign seq_loop_intf_79.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_79.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_79.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_79.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_79.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state175;
    assign seq_loop_intf_79.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state176;
    assign seq_loop_intf_79.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_79.iter_end_state1 = 452'h0;
    assign seq_loop_intf_79.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_79.one_state_loop = 1'b0;
    assign seq_loop_intf_79.one_state_block = 1'b0;
    assign seq_loop_intf_79.finish = finish;
    csv_file_dump seq_loop_csv_dumper_79;
    seq_loop_monitor #(452) seq_loop_monitor_79;
    seq_loop_intf#(452) seq_loop_intf_80(clock,reset);
    assign seq_loop_intf_80.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state176;
    assign seq_loop_intf_80.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_80.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_80.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_80.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state179;
    assign seq_loop_intf_80.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_80.post_loop_state1 = 452'h0;
    assign seq_loop_intf_80.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_80.post_loop_state2 = 452'h0;
    assign seq_loop_intf_80.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_80.post_loop_state3 = 452'h0;
    assign seq_loop_intf_80.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_80.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state178;
    assign seq_loop_intf_80.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_80.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_80.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_80.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_80.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state177;
    assign seq_loop_intf_80.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state178;
    assign seq_loop_intf_80.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_80.iter_end_state1 = 452'h0;
    assign seq_loop_intf_80.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_80.one_state_loop = 1'b0;
    assign seq_loop_intf_80.one_state_block = 1'b0;
    assign seq_loop_intf_80.finish = finish;
    csv_file_dump seq_loop_csv_dumper_80;
    seq_loop_monitor #(452) seq_loop_monitor_80;
    seq_loop_intf#(452) seq_loop_intf_81(clock,reset);
    assign seq_loop_intf_81.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state182;
    assign seq_loop_intf_81.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_81.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_81.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_81.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state185;
    assign seq_loop_intf_81.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_81.post_loop_state1 = 452'h0;
    assign seq_loop_intf_81.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_81.post_loop_state2 = 452'h0;
    assign seq_loop_intf_81.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_81.post_loop_state3 = 452'h0;
    assign seq_loop_intf_81.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_81.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state184;
    assign seq_loop_intf_81.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_81.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_81.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_81.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_81.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state183;
    assign seq_loop_intf_81.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state184;
    assign seq_loop_intf_81.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_81.iter_end_state1 = 452'h0;
    assign seq_loop_intf_81.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_81.one_state_loop = 1'b0;
    assign seq_loop_intf_81.one_state_block = 1'b0;
    assign seq_loop_intf_81.finish = finish;
    csv_file_dump seq_loop_csv_dumper_81;
    seq_loop_monitor #(452) seq_loop_monitor_81;
    seq_loop_intf#(452) seq_loop_intf_82(clock,reset);
    assign seq_loop_intf_82.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state192;
    assign seq_loop_intf_82.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_82.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_82.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_82.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state208;
    assign seq_loop_intf_82.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_82.post_loop_state1 = 452'h0;
    assign seq_loop_intf_82.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_82.post_loop_state2 = 452'h0;
    assign seq_loop_intf_82.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_82.post_loop_state3 = 452'h0;
    assign seq_loop_intf_82.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_82.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state193;
    assign seq_loop_intf_82.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_82.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_82.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_82.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_82.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state193;
    assign seq_loop_intf_82.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state207;
    assign seq_loop_intf_82.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_82.iter_end_state1 = 452'h0;
    assign seq_loop_intf_82.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_82.one_state_loop = 1'b0;
    assign seq_loop_intf_82.one_state_block = 1'b0;
    assign seq_loop_intf_82.finish = finish;
    csv_file_dump seq_loop_csv_dumper_82;
    seq_loop_monitor #(452) seq_loop_monitor_82;
    seq_loop_intf#(452) seq_loop_intf_83(clock,reset);
    assign seq_loop_intf_83.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state193;
    assign seq_loop_intf_83.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_83.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_83.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_83.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state224;
    assign seq_loop_intf_83.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_83.post_loop_state1 = 452'h0;
    assign seq_loop_intf_83.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_83.post_loop_state2 = 452'h0;
    assign seq_loop_intf_83.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_83.post_loop_state3 = 452'h0;
    assign seq_loop_intf_83.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_83.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state208;
    assign seq_loop_intf_83.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_83.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_83.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_83.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_83.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state208;
    assign seq_loop_intf_83.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state223;
    assign seq_loop_intf_83.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_83.iter_end_state1 = 452'h0;
    assign seq_loop_intf_83.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_83.one_state_loop = 1'b0;
    assign seq_loop_intf_83.one_state_block = 1'b0;
    assign seq_loop_intf_83.finish = finish;
    csv_file_dump seq_loop_csv_dumper_83;
    seq_loop_monitor #(452) seq_loop_monitor_83;
    seq_loop_intf#(452) seq_loop_intf_84(clock,reset);
    assign seq_loop_intf_84.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state208;
    assign seq_loop_intf_84.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_84.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_84.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_84.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state234;
    assign seq_loop_intf_84.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_84.post_loop_state1 = 452'h0;
    assign seq_loop_intf_84.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_84.post_loop_state2 = 452'h0;
    assign seq_loop_intf_84.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_84.post_loop_state3 = 452'h0;
    assign seq_loop_intf_84.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_84.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state224;
    assign seq_loop_intf_84.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_84.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_84.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_84.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_84.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state224;
    assign seq_loop_intf_84.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state233;
    assign seq_loop_intf_84.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_84.iter_end_state1 = 452'h0;
    assign seq_loop_intf_84.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_84.one_state_loop = 1'b0;
    assign seq_loop_intf_84.one_state_block = 1'b0;
    assign seq_loop_intf_84.finish = finish;
    csv_file_dump seq_loop_csv_dumper_84;
    seq_loop_monitor #(452) seq_loop_monitor_84;
    seq_loop_intf#(452) seq_loop_intf_85(clock,reset);
    assign seq_loop_intf_85.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state234;
    assign seq_loop_intf_85.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_85.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_85.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_85.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state240;
    assign seq_loop_intf_85.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_85.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state452;
    assign seq_loop_intf_85.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_85.post_loop_state2 = 452'h0;
    assign seq_loop_intf_85.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_85.post_loop_state3 = 452'h0;
    assign seq_loop_intf_85.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_85.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state235;
    assign seq_loop_intf_85.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_85.quit_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state236;
    assign seq_loop_intf_85.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_85.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_85.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state235;
    assign seq_loop_intf_85.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state239;
    assign seq_loop_intf_85.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_85.iter_end_state1 = 452'h0;
    assign seq_loop_intf_85.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_85.one_state_loop = 1'b0;
    assign seq_loop_intf_85.one_state_block = 1'b0;
    assign seq_loop_intf_85.finish = finish;
    csv_file_dump seq_loop_csv_dumper_85;
    seq_loop_monitor #(452) seq_loop_monitor_85;
    seq_loop_intf#(452) seq_loop_intf_86(clock,reset);
    assign seq_loop_intf_86.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state244;
    assign seq_loop_intf_86.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_86.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_86.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_86.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state249;
    assign seq_loop_intf_86.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_86.post_loop_state1 = 452'h0;
    assign seq_loop_intf_86.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_86.post_loop_state2 = 452'h0;
    assign seq_loop_intf_86.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_86.post_loop_state3 = 452'h0;
    assign seq_loop_intf_86.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_86.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state245;
    assign seq_loop_intf_86.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_86.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_86.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_86.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_86.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state245;
    assign seq_loop_intf_86.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state248;
    assign seq_loop_intf_86.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_86.iter_end_state1 = 452'h0;
    assign seq_loop_intf_86.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_86.one_state_loop = 1'b0;
    assign seq_loop_intf_86.one_state_block = 1'b0;
    assign seq_loop_intf_86.finish = finish;
    csv_file_dump seq_loop_csv_dumper_86;
    seq_loop_monitor #(452) seq_loop_monitor_86;
    seq_loop_intf#(452) seq_loop_intf_87(clock,reset);
    assign seq_loop_intf_87.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state245;
    assign seq_loop_intf_87.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_87.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_87.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_87.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state254;
    assign seq_loop_intf_87.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_87.post_loop_state1 = 452'h0;
    assign seq_loop_intf_87.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_87.post_loop_state2 = 452'h0;
    assign seq_loop_intf_87.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_87.post_loop_state3 = 452'h0;
    assign seq_loop_intf_87.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_87.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state249;
    assign seq_loop_intf_87.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_87.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_87.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_87.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_87.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state249;
    assign seq_loop_intf_87.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state253;
    assign seq_loop_intf_87.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_87.iter_end_state1 = 452'h0;
    assign seq_loop_intf_87.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_87.one_state_loop = 1'b0;
    assign seq_loop_intf_87.one_state_block = 1'b0;
    assign seq_loop_intf_87.finish = finish;
    csv_file_dump seq_loop_csv_dumper_87;
    seq_loop_monitor #(452) seq_loop_monitor_87;
    seq_loop_intf#(452) seq_loop_intf_88(clock,reset);
    assign seq_loop_intf_88.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state256;
    assign seq_loop_intf_88.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_88.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_88.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_88.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state259;
    assign seq_loop_intf_88.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_88.post_loop_state1 = 452'h0;
    assign seq_loop_intf_88.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_88.post_loop_state2 = 452'h0;
    assign seq_loop_intf_88.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_88.post_loop_state3 = 452'h0;
    assign seq_loop_intf_88.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_88.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state258;
    assign seq_loop_intf_88.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_88.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_88.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_88.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_88.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state257;
    assign seq_loop_intf_88.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state258;
    assign seq_loop_intf_88.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_88.iter_end_state1 = 452'h0;
    assign seq_loop_intf_88.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_88.one_state_loop = 1'b0;
    assign seq_loop_intf_88.one_state_block = 1'b0;
    assign seq_loop_intf_88.finish = finish;
    csv_file_dump seq_loop_csv_dumper_88;
    seq_loop_monitor #(452) seq_loop_monitor_88;
    seq_loop_intf#(452) seq_loop_intf_89(clock,reset);
    assign seq_loop_intf_89.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state258;
    assign seq_loop_intf_89.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_89.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_89.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_89.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state452;
    assign seq_loop_intf_89.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_89.post_loop_state1 = 452'h0;
    assign seq_loop_intf_89.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_89.post_loop_state2 = 452'h0;
    assign seq_loop_intf_89.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_89.post_loop_state3 = 452'h0;
    assign seq_loop_intf_89.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_89.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state259;
    assign seq_loop_intf_89.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_89.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_89.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_89.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_89.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state259;
    assign seq_loop_intf_89.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state264;
    assign seq_loop_intf_89.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_89.iter_end_state1 = 452'h0;
    assign seq_loop_intf_89.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_89.one_state_loop = 1'b0;
    assign seq_loop_intf_89.one_state_block = 1'b0;
    assign seq_loop_intf_89.finish = finish;
    csv_file_dump seq_loop_csv_dumper_89;
    seq_loop_monitor #(452) seq_loop_monitor_89;
    seq_loop_intf#(452) seq_loop_intf_90(clock,reset);
    assign seq_loop_intf_90.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state2;
    assign seq_loop_intf_90.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_90.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_90.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_90.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state5;
    assign seq_loop_intf_90.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_90.post_loop_state1 = 452'h0;
    assign seq_loop_intf_90.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_90.post_loop_state2 = 452'h0;
    assign seq_loop_intf_90.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_90.post_loop_state3 = 452'h0;
    assign seq_loop_intf_90.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_90.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state3;
    assign seq_loop_intf_90.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_90.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_90.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_90.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_90.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state3;
    assign seq_loop_intf_90.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state4;
    assign seq_loop_intf_90.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_90.iter_end_state1 = 452'h0;
    assign seq_loop_intf_90.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_90.one_state_loop = 1'b0;
    assign seq_loop_intf_90.one_state_block = 1'b0;
    assign seq_loop_intf_90.finish = finish;
    csv_file_dump seq_loop_csv_dumper_90;
    seq_loop_monitor #(452) seq_loop_monitor_90;
    seq_loop_intf#(452) seq_loop_intf_91(clock,reset);
    assign seq_loop_intf_91.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state7;
    assign seq_loop_intf_91.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_91.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_91.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_91.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state10;
    assign seq_loop_intf_91.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_91.post_loop_state1 = 452'h0;
    assign seq_loop_intf_91.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_91.post_loop_state2 = 452'h0;
    assign seq_loop_intf_91.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_91.post_loop_state3 = 452'h0;
    assign seq_loop_intf_91.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_91.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state8;
    assign seq_loop_intf_91.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_91.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_91.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_91.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_91.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state8;
    assign seq_loop_intf_91.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state9;
    assign seq_loop_intf_91.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_91.iter_end_state1 = 452'h0;
    assign seq_loop_intf_91.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_91.one_state_loop = 1'b0;
    assign seq_loop_intf_91.one_state_block = 1'b0;
    assign seq_loop_intf_91.finish = finish;
    csv_file_dump seq_loop_csv_dumper_91;
    seq_loop_monitor #(452) seq_loop_monitor_91;
    seq_loop_intf#(452) seq_loop_intf_92(clock,reset);
    assign seq_loop_intf_92.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state12;
    assign seq_loop_intf_92.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_92.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_92.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_92.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state19;
    assign seq_loop_intf_92.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_92.post_loop_state1 = 452'h0;
    assign seq_loop_intf_92.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_92.post_loop_state2 = 452'h0;
    assign seq_loop_intf_92.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_92.post_loop_state3 = 452'h0;
    assign seq_loop_intf_92.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_92.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state13;
    assign seq_loop_intf_92.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_92.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_92.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_92.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_92.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state13;
    assign seq_loop_intf_92.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state18;
    assign seq_loop_intf_92.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_92.iter_end_state1 = 452'h0;
    assign seq_loop_intf_92.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_92.one_state_loop = 1'b0;
    assign seq_loop_intf_92.one_state_block = 1'b0;
    assign seq_loop_intf_92.finish = finish;
    csv_file_dump seq_loop_csv_dumper_92;
    seq_loop_monitor #(452) seq_loop_monitor_92;
    seq_loop_intf#(452) seq_loop_intf_93(clock,reset);
    assign seq_loop_intf_93.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state21;
    assign seq_loop_intf_93.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_93.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_93.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_93.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state24;
    assign seq_loop_intf_93.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_93.post_loop_state1 = 452'h0;
    assign seq_loop_intf_93.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_93.post_loop_state2 = 452'h0;
    assign seq_loop_intf_93.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_93.post_loop_state3 = 452'h0;
    assign seq_loop_intf_93.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_93.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state23;
    assign seq_loop_intf_93.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_93.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_93.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_93.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_93.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state22;
    assign seq_loop_intf_93.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state23;
    assign seq_loop_intf_93.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_93.iter_end_state1 = 452'h0;
    assign seq_loop_intf_93.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_93.one_state_loop = 1'b0;
    assign seq_loop_intf_93.one_state_block = 1'b0;
    assign seq_loop_intf_93.finish = finish;
    csv_file_dump seq_loop_csv_dumper_93;
    seq_loop_monitor #(452) seq_loop_monitor_93;
    seq_loop_intf#(452) seq_loop_intf_94(clock,reset);
    assign seq_loop_intf_94.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state30;
    assign seq_loop_intf_94.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_94.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_94.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_94.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state34;
    assign seq_loop_intf_94.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_94.post_loop_state1 = 452'h0;
    assign seq_loop_intf_94.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_94.post_loop_state2 = 452'h0;
    assign seq_loop_intf_94.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_94.post_loop_state3 = 452'h0;
    assign seq_loop_intf_94.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_94.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state31;
    assign seq_loop_intf_94.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_94.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_94.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_94.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_94.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state31;
    assign seq_loop_intf_94.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state33;
    assign seq_loop_intf_94.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_94.iter_end_state1 = 452'h0;
    assign seq_loop_intf_94.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_94.one_state_loop = 1'b0;
    assign seq_loop_intf_94.one_state_block = 1'b0;
    assign seq_loop_intf_94.finish = finish;
    csv_file_dump seq_loop_csv_dumper_94;
    seq_loop_monitor #(452) seq_loop_monitor_94;
    seq_loop_intf#(452) seq_loop_intf_95(clock,reset);
    assign seq_loop_intf_95.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state36;
    assign seq_loop_intf_95.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_95.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_95.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_95.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state40;
    assign seq_loop_intf_95.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_95.post_loop_state1 = 452'h0;
    assign seq_loop_intf_95.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_95.post_loop_state2 = 452'h0;
    assign seq_loop_intf_95.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_95.post_loop_state3 = 452'h0;
    assign seq_loop_intf_95.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_95.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state37;
    assign seq_loop_intf_95.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_95.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_95.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_95.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_95.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state37;
    assign seq_loop_intf_95.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state39;
    assign seq_loop_intf_95.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_95.iter_end_state1 = 452'h0;
    assign seq_loop_intf_95.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_95.one_state_loop = 1'b0;
    assign seq_loop_intf_95.one_state_block = 1'b0;
    assign seq_loop_intf_95.finish = finish;
    csv_file_dump seq_loop_csv_dumper_95;
    seq_loop_monitor #(452) seq_loop_monitor_95;
    seq_loop_intf#(452) seq_loop_intf_96(clock,reset);
    assign seq_loop_intf_96.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state40;
    assign seq_loop_intf_96.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_96.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_96.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_96.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state44;
    assign seq_loop_intf_96.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_96.post_loop_state1 = 452'h0;
    assign seq_loop_intf_96.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_96.post_loop_state2 = 452'h0;
    assign seq_loop_intf_96.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_96.post_loop_state3 = 452'h0;
    assign seq_loop_intf_96.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_96.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state41;
    assign seq_loop_intf_96.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_96.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_96.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_96.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_96.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state41;
    assign seq_loop_intf_96.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state43;
    assign seq_loop_intf_96.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_96.iter_end_state1 = 452'h0;
    assign seq_loop_intf_96.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_96.one_state_loop = 1'b0;
    assign seq_loop_intf_96.one_state_block = 1'b0;
    assign seq_loop_intf_96.finish = finish;
    csv_file_dump seq_loop_csv_dumper_96;
    seq_loop_monitor #(452) seq_loop_monitor_96;
    seq_loop_intf#(452) seq_loop_intf_97(clock,reset);
    assign seq_loop_intf_97.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state46;
    assign seq_loop_intf_97.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_97.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_97.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_97.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state51;
    assign seq_loop_intf_97.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_97.post_loop_state1 = 452'h0;
    assign seq_loop_intf_97.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_97.post_loop_state2 = 452'h0;
    assign seq_loop_intf_97.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_97.post_loop_state3 = 452'h0;
    assign seq_loop_intf_97.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_97.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state47;
    assign seq_loop_intf_97.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_97.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_97.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_97.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_97.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state47;
    assign seq_loop_intf_97.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state50;
    assign seq_loop_intf_97.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_97.iter_end_state1 = 452'h0;
    assign seq_loop_intf_97.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_97.one_state_loop = 1'b0;
    assign seq_loop_intf_97.one_state_block = 1'b0;
    assign seq_loop_intf_97.finish = finish;
    csv_file_dump seq_loop_csv_dumper_97;
    seq_loop_monitor #(452) seq_loop_monitor_97;
    seq_loop_intf#(452) seq_loop_intf_98(clock,reset);
    assign seq_loop_intf_98.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state55;
    assign seq_loop_intf_98.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_98.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_98.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_98.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state58;
    assign seq_loop_intf_98.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_98.post_loop_state1 = 452'h0;
    assign seq_loop_intf_98.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_98.post_loop_state2 = 452'h0;
    assign seq_loop_intf_98.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_98.post_loop_state3 = 452'h0;
    assign seq_loop_intf_98.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_98.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state56;
    assign seq_loop_intf_98.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_98.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_98.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_98.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_98.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state56;
    assign seq_loop_intf_98.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state57;
    assign seq_loop_intf_98.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_98.iter_end_state1 = 452'h0;
    assign seq_loop_intf_98.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_98.one_state_loop = 1'b0;
    assign seq_loop_intf_98.one_state_block = 1'b0;
    assign seq_loop_intf_98.finish = finish;
    csv_file_dump seq_loop_csv_dumper_98;
    seq_loop_monitor #(452) seq_loop_monitor_98;
    seq_loop_intf#(452) seq_loop_intf_99(clock,reset);
    assign seq_loop_intf_99.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state56;
    assign seq_loop_intf_99.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_99.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_99.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_99.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state62;
    assign seq_loop_intf_99.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_99.post_loop_state1 = 452'h0;
    assign seq_loop_intf_99.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_99.post_loop_state2 = 452'h0;
    assign seq_loop_intf_99.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_99.post_loop_state3 = 452'h0;
    assign seq_loop_intf_99.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_99.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state58;
    assign seq_loop_intf_99.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_99.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_99.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_99.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_99.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state58;
    assign seq_loop_intf_99.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state61;
    assign seq_loop_intf_99.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_99.iter_end_state1 = 452'h0;
    assign seq_loop_intf_99.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_99.one_state_loop = 1'b0;
    assign seq_loop_intf_99.one_state_block = 1'b0;
    assign seq_loop_intf_99.finish = finish;
    csv_file_dump seq_loop_csv_dumper_99;
    seq_loop_monitor #(452) seq_loop_monitor_99;
    seq_loop_intf#(452) seq_loop_intf_100(clock,reset);
    assign seq_loop_intf_100.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state62;
    assign seq_loop_intf_100.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_100.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_100.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_100.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state65;
    assign seq_loop_intf_100.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_100.post_loop_state1 = 452'h0;
    assign seq_loop_intf_100.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_100.post_loop_state2 = 452'h0;
    assign seq_loop_intf_100.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_100.post_loop_state3 = 452'h0;
    assign seq_loop_intf_100.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_100.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state64;
    assign seq_loop_intf_100.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_100.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_100.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_100.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_100.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state63;
    assign seq_loop_intf_100.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state64;
    assign seq_loop_intf_100.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_100.iter_end_state1 = 452'h0;
    assign seq_loop_intf_100.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_100.one_state_loop = 1'b0;
    assign seq_loop_intf_100.one_state_block = 1'b0;
    assign seq_loop_intf_100.finish = finish;
    csv_file_dump seq_loop_csv_dumper_100;
    seq_loop_monitor #(452) seq_loop_monitor_100;
    seq_loop_intf#(452) seq_loop_intf_101(clock,reset);
    assign seq_loop_intf_101.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state64;
    assign seq_loop_intf_101.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_101.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_101.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_101.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state69;
    assign seq_loop_intf_101.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_101.post_loop_state1 = 452'h0;
    assign seq_loop_intf_101.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_101.post_loop_state2 = 452'h0;
    assign seq_loop_intf_101.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_101.post_loop_state3 = 452'h0;
    assign seq_loop_intf_101.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_101.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state65;
    assign seq_loop_intf_101.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_101.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_101.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_101.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_101.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state65;
    assign seq_loop_intf_101.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state68;
    assign seq_loop_intf_101.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_101.iter_end_state1 = 452'h0;
    assign seq_loop_intf_101.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_101.one_state_loop = 1'b0;
    assign seq_loop_intf_101.one_state_block = 1'b0;
    assign seq_loop_intf_101.finish = finish;
    csv_file_dump seq_loop_csv_dumper_101;
    seq_loop_monitor #(452) seq_loop_monitor_101;
    seq_loop_intf#(452) seq_loop_intf_102(clock,reset);
    assign seq_loop_intf_102.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state69;
    assign seq_loop_intf_102.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_102.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_102.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_102.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state85;
    assign seq_loop_intf_102.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_102.post_loop_state1 = 452'h0;
    assign seq_loop_intf_102.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_102.post_loop_state2 = 452'h0;
    assign seq_loop_intf_102.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_102.post_loop_state3 = 452'h0;
    assign seq_loop_intf_102.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_102.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state70;
    assign seq_loop_intf_102.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_102.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_102.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_102.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_102.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state70;
    assign seq_loop_intf_102.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state84;
    assign seq_loop_intf_102.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_102.iter_end_state1 = 452'h0;
    assign seq_loop_intf_102.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_102.one_state_loop = 1'b0;
    assign seq_loop_intf_102.one_state_block = 1'b0;
    assign seq_loop_intf_102.finish = finish;
    csv_file_dump seq_loop_csv_dumper_102;
    seq_loop_monitor #(452) seq_loop_monitor_102;
    seq_loop_intf#(452) seq_loop_intf_103(clock,reset);
    assign seq_loop_intf_103.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state85;
    assign seq_loop_intf_103.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_103.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_103.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_103.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state89;
    assign seq_loop_intf_103.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_103.post_loop_state1 = 452'h0;
    assign seq_loop_intf_103.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_103.post_loop_state2 = 452'h0;
    assign seq_loop_intf_103.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_103.post_loop_state3 = 452'h0;
    assign seq_loop_intf_103.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_103.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state86;
    assign seq_loop_intf_103.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_103.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_103.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_103.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_103.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state86;
    assign seq_loop_intf_103.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state88;
    assign seq_loop_intf_103.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_103.iter_end_state1 = 452'h0;
    assign seq_loop_intf_103.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_103.one_state_loop = 1'b0;
    assign seq_loop_intf_103.one_state_block = 1'b0;
    assign seq_loop_intf_103.finish = finish;
    csv_file_dump seq_loop_csv_dumper_103;
    seq_loop_monitor #(452) seq_loop_monitor_103;
    seq_loop_intf#(452) seq_loop_intf_104(clock,reset);
    assign seq_loop_intf_104.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state89;
    assign seq_loop_intf_104.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_104.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_104.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_104.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state92;
    assign seq_loop_intf_104.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_104.post_loop_state1 = 452'h0;
    assign seq_loop_intf_104.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_104.post_loop_state2 = 452'h0;
    assign seq_loop_intf_104.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_104.post_loop_state3 = 452'h0;
    assign seq_loop_intf_104.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_104.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state90;
    assign seq_loop_intf_104.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_104.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_104.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_104.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_104.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state90;
    assign seq_loop_intf_104.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state91;
    assign seq_loop_intf_104.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_104.iter_end_state1 = 452'h0;
    assign seq_loop_intf_104.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_104.one_state_loop = 1'b0;
    assign seq_loop_intf_104.one_state_block = 1'b0;
    assign seq_loop_intf_104.finish = finish;
    csv_file_dump seq_loop_csv_dumper_104;
    seq_loop_monitor #(452) seq_loop_monitor_104;
    seq_loop_intf#(452) seq_loop_intf_105(clock,reset);
    assign seq_loop_intf_105.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state96;
    assign seq_loop_intf_105.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_105.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_105.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_105.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state101;
    assign seq_loop_intf_105.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_105.post_loop_state1 = 452'h0;
    assign seq_loop_intf_105.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_105.post_loop_state2 = 452'h0;
    assign seq_loop_intf_105.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_105.post_loop_state3 = 452'h0;
    assign seq_loop_intf_105.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_105.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state97;
    assign seq_loop_intf_105.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_105.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_105.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_105.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_105.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state97;
    assign seq_loop_intf_105.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state100;
    assign seq_loop_intf_105.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_105.iter_end_state1 = 452'h0;
    assign seq_loop_intf_105.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_105.one_state_loop = 1'b0;
    assign seq_loop_intf_105.one_state_block = 1'b0;
    assign seq_loop_intf_105.finish = finish;
    csv_file_dump seq_loop_csv_dumper_105;
    seq_loop_monitor #(452) seq_loop_monitor_105;
    seq_loop_intf#(452) seq_loop_intf_106(clock,reset);
    assign seq_loop_intf_106.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state103;
    assign seq_loop_intf_106.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_106.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_106.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_106.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state452;
    assign seq_loop_intf_106.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_106.post_loop_state1 = 452'h0;
    assign seq_loop_intf_106.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_106.post_loop_state2 = 452'h0;
    assign seq_loop_intf_106.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_106.post_loop_state3 = 452'h0;
    assign seq_loop_intf_106.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_106.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state104;
    assign seq_loop_intf_106.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_106.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_106.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_106.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_106.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state104;
    assign seq_loop_intf_106.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state105;
    assign seq_loop_intf_106.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_106.iter_end_state1 = 452'h0;
    assign seq_loop_intf_106.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_106.one_state_loop = 1'b0;
    assign seq_loop_intf_106.one_state_block = 1'b0;
    assign seq_loop_intf_106.finish = finish;
    csv_file_dump seq_loop_csv_dumper_106;
    seq_loop_monitor #(452) seq_loop_monitor_106;
    seq_loop_intf#(452) seq_loop_intf_107(clock,reset);
    assign seq_loop_intf_107.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state275;
    assign seq_loop_intf_107.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_107.pre_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state276;
    assign seq_loop_intf_107.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_107.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state276;
    assign seq_loop_intf_107.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_107.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state280;
    assign seq_loop_intf_107.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_107.post_loop_state2 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state279;
    assign seq_loop_intf_107.post_states_valid[2] = 1'b1;
    assign seq_loop_intf_107.post_loop_state3 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state281;
    assign seq_loop_intf_107.post_states_valid[3] = 1'b1;
    assign seq_loop_intf_107.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state277;
    assign seq_loop_intf_107.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_107.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_107.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_107.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_107.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state277;
    assign seq_loop_intf_107.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state278;
    assign seq_loop_intf_107.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_107.iter_end_state1 = 452'h0;
    assign seq_loop_intf_107.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_107.one_state_loop = 1'b0;
    assign seq_loop_intf_107.one_state_block = 1'b0;
    assign seq_loop_intf_107.finish = finish;
    csv_file_dump seq_loop_csv_dumper_107;
    seq_loop_monitor #(452) seq_loop_monitor_107;
    seq_loop_intf#(452) seq_loop_intf_108(clock,reset);
    assign seq_loop_intf_108.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state275;
    assign seq_loop_intf_108.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_108.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_108.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_108.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state278;
    assign seq_loop_intf_108.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_108.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state280;
    assign seq_loop_intf_108.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_108.post_loop_state2 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state279;
    assign seq_loop_intf_108.post_states_valid[2] = 1'b1;
    assign seq_loop_intf_108.post_loop_state3 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state281;
    assign seq_loop_intf_108.post_states_valid[3] = 1'b1;
    assign seq_loop_intf_108.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state277;
    assign seq_loop_intf_108.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_108.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_108.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_108.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_108.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state276;
    assign seq_loop_intf_108.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state277;
    assign seq_loop_intf_108.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_108.iter_end_state1 = 452'h0;
    assign seq_loop_intf_108.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_108.one_state_loop = 1'b0;
    assign seq_loop_intf_108.one_state_block = 1'b0;
    assign seq_loop_intf_108.finish = finish;
    csv_file_dump seq_loop_csv_dumper_108;
    seq_loop_monitor #(452) seq_loop_monitor_108;
    seq_loop_intf#(452) seq_loop_intf_109(clock,reset);
    assign seq_loop_intf_109.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state277;
    assign seq_loop_intf_109.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_109.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_109.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_109.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state281;
    assign seq_loop_intf_109.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_109.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state282;
    assign seq_loop_intf_109.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_109.post_loop_state2 = 452'h0;
    assign seq_loop_intf_109.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_109.post_loop_state3 = 452'h0;
    assign seq_loop_intf_109.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_109.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state280;
    assign seq_loop_intf_109.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_109.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_109.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_109.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_109.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state279;
    assign seq_loop_intf_109.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state280;
    assign seq_loop_intf_109.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_109.iter_end_state1 = 452'h0;
    assign seq_loop_intf_109.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_109.one_state_loop = 1'b0;
    assign seq_loop_intf_109.one_state_block = 1'b0;
    assign seq_loop_intf_109.finish = finish;
    csv_file_dump seq_loop_csv_dumper_109;
    seq_loop_monitor #(452) seq_loop_monitor_109;
    seq_loop_intf#(452) seq_loop_intf_110(clock,reset);
    assign seq_loop_intf_110.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state277;
    assign seq_loop_intf_110.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_110.pre_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state279;
    assign seq_loop_intf_110.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_110.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state279;
    assign seq_loop_intf_110.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_110.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state282;
    assign seq_loop_intf_110.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_110.post_loop_state2 = 452'h0;
    assign seq_loop_intf_110.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_110.post_loop_state3 = 452'h0;
    assign seq_loop_intf_110.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_110.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state280;
    assign seq_loop_intf_110.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_110.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_110.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_110.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_110.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state280;
    assign seq_loop_intf_110.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state281;
    assign seq_loop_intf_110.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_110.iter_end_state1 = 452'h0;
    assign seq_loop_intf_110.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_110.one_state_loop = 1'b0;
    assign seq_loop_intf_110.one_state_block = 1'b0;
    assign seq_loop_intf_110.finish = finish;
    csv_file_dump seq_loop_csv_dumper_110;
    seq_loop_monitor #(452) seq_loop_monitor_110;
    seq_loop_intf#(452) seq_loop_intf_111(clock,reset);
    assign seq_loop_intf_111.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state286;
    assign seq_loop_intf_111.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_111.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_111.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_111.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state289;
    assign seq_loop_intf_111.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_111.post_loop_state1 = 452'h0;
    assign seq_loop_intf_111.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_111.post_loop_state2 = 452'h0;
    assign seq_loop_intf_111.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_111.post_loop_state3 = 452'h0;
    assign seq_loop_intf_111.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_111.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state287;
    assign seq_loop_intf_111.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_111.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_111.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_111.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_111.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state287;
    assign seq_loop_intf_111.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state288;
    assign seq_loop_intf_111.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_111.iter_end_state1 = 452'h0;
    assign seq_loop_intf_111.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_111.one_state_loop = 1'b0;
    assign seq_loop_intf_111.one_state_block = 1'b0;
    assign seq_loop_intf_111.finish = finish;
    csv_file_dump seq_loop_csv_dumper_111;
    seq_loop_monitor #(452) seq_loop_monitor_111;
    seq_loop_intf#(452) seq_loop_intf_112(clock,reset);
    assign seq_loop_intf_112.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state287;
    assign seq_loop_intf_112.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_112.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_112.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_112.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state282;
    assign seq_loop_intf_112.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_112.post_loop_state1 = 452'h0;
    assign seq_loop_intf_112.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_112.post_loop_state2 = 452'h0;
    assign seq_loop_intf_112.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_112.post_loop_state3 = 452'h0;
    assign seq_loop_intf_112.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_112.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state289;
    assign seq_loop_intf_112.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_112.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_112.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_112.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_112.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state289;
    assign seq_loop_intf_112.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state294;
    assign seq_loop_intf_112.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_112.iter_end_state1 = 452'h0;
    assign seq_loop_intf_112.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_112.one_state_loop = 1'b0;
    assign seq_loop_intf_112.one_state_block = 1'b0;
    assign seq_loop_intf_112.finish = finish;
    csv_file_dump seq_loop_csv_dumper_112;
    seq_loop_monitor #(452) seq_loop_monitor_112;
    seq_loop_intf#(452) seq_loop_intf_113(clock,reset);
    assign seq_loop_intf_113.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state280;
    assign seq_loop_intf_113.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_113.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_113.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_113.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state295;
    assign seq_loop_intf_113.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_113.post_loop_state1 = 452'h0;
    assign seq_loop_intf_113.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_113.post_loop_state2 = 452'h0;
    assign seq_loop_intf_113.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_113.post_loop_state3 = 452'h0;
    assign seq_loop_intf_113.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_113.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state282;
    assign seq_loop_intf_113.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_113.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_113.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_113.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_113.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state282;
    assign seq_loop_intf_113.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state289;
    assign seq_loop_intf_113.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_113.iter_end_state1 = 452'h0;
    assign seq_loop_intf_113.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_113.one_state_loop = 1'b0;
    assign seq_loop_intf_113.one_state_block = 1'b0;
    assign seq_loop_intf_113.finish = finish;
    csv_file_dump seq_loop_csv_dumper_113;
    seq_loop_monitor #(452) seq_loop_monitor_113;
    seq_loop_intf#(452) seq_loop_intf_114(clock,reset);
    assign seq_loop_intf_114.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state304;
    assign seq_loop_intf_114.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_114.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_114.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_114.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state320;
    assign seq_loop_intf_114.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_114.post_loop_state1 = 452'h0;
    assign seq_loop_intf_114.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_114.post_loop_state2 = 452'h0;
    assign seq_loop_intf_114.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_114.post_loop_state3 = 452'h0;
    assign seq_loop_intf_114.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_114.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state316;
    assign seq_loop_intf_114.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_114.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_114.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_114.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_114.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state316;
    assign seq_loop_intf_114.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state319;
    assign seq_loop_intf_114.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_114.iter_end_state1 = 452'h0;
    assign seq_loop_intf_114.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_114.one_state_loop = 1'b0;
    assign seq_loop_intf_114.one_state_block = 1'b0;
    assign seq_loop_intf_114.finish = finish;
    csv_file_dump seq_loop_csv_dumper_114;
    seq_loop_monitor #(452) seq_loop_monitor_114;
    seq_loop_intf#(452) seq_loop_intf_115(clock,reset);
    assign seq_loop_intf_115.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state304;
    assign seq_loop_intf_115.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_115.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_115.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_115.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state307;
    assign seq_loop_intf_115.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_115.post_loop_state1 = 452'h0;
    assign seq_loop_intf_115.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_115.post_loop_state2 = 452'h0;
    assign seq_loop_intf_115.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_115.post_loop_state3 = 452'h0;
    assign seq_loop_intf_115.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_115.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state305;
    assign seq_loop_intf_115.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_115.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_115.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_115.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_115.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state305;
    assign seq_loop_intf_115.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state306;
    assign seq_loop_intf_115.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_115.iter_end_state1 = 452'h0;
    assign seq_loop_intf_115.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_115.one_state_loop = 1'b0;
    assign seq_loop_intf_115.one_state_block = 1'b0;
    assign seq_loop_intf_115.finish = finish;
    csv_file_dump seq_loop_csv_dumper_115;
    seq_loop_monitor #(452) seq_loop_monitor_115;
    seq_loop_intf#(452) seq_loop_intf_116(clock,reset);
    assign seq_loop_intf_116.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state305;
    assign seq_loop_intf_116.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_116.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_116.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_116.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state313;
    assign seq_loop_intf_116.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_116.post_loop_state1 = 452'h0;
    assign seq_loop_intf_116.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_116.post_loop_state2 = 452'h0;
    assign seq_loop_intf_116.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_116.post_loop_state3 = 452'h0;
    assign seq_loop_intf_116.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_116.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state307;
    assign seq_loop_intf_116.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_116.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_116.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_116.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_116.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state307;
    assign seq_loop_intf_116.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state312;
    assign seq_loop_intf_116.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_116.iter_end_state1 = 452'h0;
    assign seq_loop_intf_116.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_116.one_state_loop = 1'b0;
    assign seq_loop_intf_116.one_state_block = 1'b0;
    assign seq_loop_intf_116.finish = finish;
    csv_file_dump seq_loop_csv_dumper_116;
    seq_loop_monitor #(452) seq_loop_monitor_116;
    seq_loop_intf#(452) seq_loop_intf_117(clock,reset);
    assign seq_loop_intf_117.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state315;
    assign seq_loop_intf_117.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_117.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_117.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_117.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state327;
    assign seq_loop_intf_117.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_117.post_loop_state1 = 452'h0;
    assign seq_loop_intf_117.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_117.post_loop_state2 = 452'h0;
    assign seq_loop_intf_117.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_117.post_loop_state3 = 452'h0;
    assign seq_loop_intf_117.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_117.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state323;
    assign seq_loop_intf_117.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_117.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_117.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_117.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_117.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state323;
    assign seq_loop_intf_117.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state326;
    assign seq_loop_intf_117.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_117.iter_end_state1 = 452'h0;
    assign seq_loop_intf_117.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_117.one_state_loop = 1'b0;
    assign seq_loop_intf_117.one_state_block = 1'b0;
    assign seq_loop_intf_117.finish = finish;
    csv_file_dump seq_loop_csv_dumper_117;
    seq_loop_monitor #(452) seq_loop_monitor_117;
    seq_loop_intf#(452) seq_loop_intf_118(clock,reset);
    assign seq_loop_intf_118.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state329;
    assign seq_loop_intf_118.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_118.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_118.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_118.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state337;
    assign seq_loop_intf_118.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_118.post_loop_state1 = 452'h0;
    assign seq_loop_intf_118.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_118.post_loop_state2 = 452'h0;
    assign seq_loop_intf_118.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_118.post_loop_state3 = 452'h0;
    assign seq_loop_intf_118.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_118.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state330;
    assign seq_loop_intf_118.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_118.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_118.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_118.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_118.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state330;
    assign seq_loop_intf_118.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state336;
    assign seq_loop_intf_118.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_118.iter_end_state1 = 452'h0;
    assign seq_loop_intf_118.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_118.one_state_loop = 1'b0;
    assign seq_loop_intf_118.one_state_block = 1'b0;
    assign seq_loop_intf_118.finish = finish;
    csv_file_dump seq_loop_csv_dumper_118;
    seq_loop_monitor #(452) seq_loop_monitor_118;
    seq_loop_intf#(452) seq_loop_intf_119(clock,reset);
    assign seq_loop_intf_119.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state282;
    assign seq_loop_intf_119.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_119.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_119.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_119.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state340;
    assign seq_loop_intf_119.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_119.post_loop_state1 = 452'h0;
    assign seq_loop_intf_119.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_119.post_loop_state2 = 452'h0;
    assign seq_loop_intf_119.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_119.post_loop_state3 = 452'h0;
    assign seq_loop_intf_119.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_119.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state295;
    assign seq_loop_intf_119.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_119.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_119.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_119.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_119.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state295;
    assign seq_loop_intf_119.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state339;
    assign seq_loop_intf_119.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_119.iter_end_state1 = 452'h0;
    assign seq_loop_intf_119.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_119.one_state_loop = 1'b0;
    assign seq_loop_intf_119.one_state_block = 1'b0;
    assign seq_loop_intf_119.finish = finish;
    csv_file_dump seq_loop_csv_dumper_119;
    seq_loop_monitor #(452) seq_loop_monitor_119;
    seq_loop_intf#(452) seq_loop_intf_120(clock,reset);
    assign seq_loop_intf_120.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state350;
    assign seq_loop_intf_120.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_120.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_120.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_120.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state368;
    assign seq_loop_intf_120.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_120.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state366;
    assign seq_loop_intf_120.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_120.post_loop_state2 = 452'h0;
    assign seq_loop_intf_120.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_120.post_loop_state3 = 452'h0;
    assign seq_loop_intf_120.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_120.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state351;
    assign seq_loop_intf_120.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_120.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_120.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_120.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_120.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state351;
    assign seq_loop_intf_120.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state365;
    assign seq_loop_intf_120.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_120.iter_end_state1 = 452'h0;
    assign seq_loop_intf_120.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_120.one_state_loop = 1'b0;
    assign seq_loop_intf_120.one_state_block = 1'b0;
    assign seq_loop_intf_120.finish = finish;
    csv_file_dump seq_loop_csv_dumper_120;
    seq_loop_monitor #(452) seq_loop_monitor_120;
    seq_loop_intf#(452) seq_loop_intf_121(clock,reset);
    assign seq_loop_intf_121.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state351;
    assign seq_loop_intf_121.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_121.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_121.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_121.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state368;
    assign seq_loop_intf_121.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_121.post_loop_state1 = 452'h0;
    assign seq_loop_intf_121.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_121.post_loop_state2 = 452'h0;
    assign seq_loop_intf_121.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_121.post_loop_state3 = 452'h0;
    assign seq_loop_intf_121.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_121.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state366;
    assign seq_loop_intf_121.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_121.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_121.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_121.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_121.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state366;
    assign seq_loop_intf_121.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state367;
    assign seq_loop_intf_121.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_121.iter_end_state1 = 452'h0;
    assign seq_loop_intf_121.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_121.one_state_loop = 1'b0;
    assign seq_loop_intf_121.one_state_block = 1'b0;
    assign seq_loop_intf_121.finish = finish;
    csv_file_dump seq_loop_csv_dumper_121;
    seq_loop_monitor #(452) seq_loop_monitor_121;
    seq_loop_intf#(452) seq_loop_intf_122(clock,reset);
    assign seq_loop_intf_122.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state351;
    assign seq_loop_intf_122.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_122.pre_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state366;
    assign seq_loop_intf_122.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_122.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state370;
    assign seq_loop_intf_122.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_122.post_loop_state1 = 452'h0;
    assign seq_loop_intf_122.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_122.post_loop_state2 = 452'h0;
    assign seq_loop_intf_122.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_122.post_loop_state3 = 452'h0;
    assign seq_loop_intf_122.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_122.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state368;
    assign seq_loop_intf_122.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_122.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_122.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_122.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_122.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state368;
    assign seq_loop_intf_122.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state369;
    assign seq_loop_intf_122.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_122.iter_end_state1 = 452'h0;
    assign seq_loop_intf_122.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_122.one_state_loop = 1'b0;
    assign seq_loop_intf_122.one_state_block = 1'b0;
    assign seq_loop_intf_122.finish = finish;
    csv_file_dump seq_loop_csv_dumper_122;
    seq_loop_monitor #(452) seq_loop_monitor_122;
    seq_loop_intf#(452) seq_loop_intf_123(clock,reset);
    assign seq_loop_intf_123.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state381;
    assign seq_loop_intf_123.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_123.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_123.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_123.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state386;
    assign seq_loop_intf_123.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_123.post_loop_state1 = 452'h0;
    assign seq_loop_intf_123.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_123.post_loop_state2 = 452'h0;
    assign seq_loop_intf_123.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_123.post_loop_state3 = 452'h0;
    assign seq_loop_intf_123.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_123.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state382;
    assign seq_loop_intf_123.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_123.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_123.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_123.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_123.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state382;
    assign seq_loop_intf_123.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state385;
    assign seq_loop_intf_123.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_123.iter_end_state1 = 452'h0;
    assign seq_loop_intf_123.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_123.one_state_loop = 1'b0;
    assign seq_loop_intf_123.one_state_block = 1'b0;
    assign seq_loop_intf_123.finish = finish;
    csv_file_dump seq_loop_csv_dumper_123;
    seq_loop_monitor #(452) seq_loop_monitor_123;
    seq_loop_intf#(452) seq_loop_intf_124(clock,reset);
    assign seq_loop_intf_124.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state382;
    assign seq_loop_intf_124.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_124.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_124.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_124.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state394;
    assign seq_loop_intf_124.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_124.post_loop_state1 = 452'h0;
    assign seq_loop_intf_124.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_124.post_loop_state2 = 452'h0;
    assign seq_loop_intf_124.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_124.post_loop_state3 = 452'h0;
    assign seq_loop_intf_124.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_124.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state386;
    assign seq_loop_intf_124.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_124.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_124.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_124.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_124.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state386;
    assign seq_loop_intf_124.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state393;
    assign seq_loop_intf_124.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_124.iter_end_state1 = 452'h0;
    assign seq_loop_intf_124.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_124.one_state_loop = 1'b0;
    assign seq_loop_intf_124.one_state_block = 1'b0;
    assign seq_loop_intf_124.finish = finish;
    csv_file_dump seq_loop_csv_dumper_124;
    seq_loop_monitor #(452) seq_loop_monitor_124;
    seq_loop_intf#(452) seq_loop_intf_125(clock,reset);
    assign seq_loop_intf_125.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state394;
    assign seq_loop_intf_125.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_125.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_125.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_125.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state398;
    assign seq_loop_intf_125.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_125.post_loop_state1 = 452'h0;
    assign seq_loop_intf_125.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_125.post_loop_state2 = 452'h0;
    assign seq_loop_intf_125.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_125.post_loop_state3 = 452'h0;
    assign seq_loop_intf_125.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_125.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state395;
    assign seq_loop_intf_125.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_125.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_125.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_125.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_125.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state395;
    assign seq_loop_intf_125.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state397;
    assign seq_loop_intf_125.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_125.iter_end_state1 = 452'h0;
    assign seq_loop_intf_125.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_125.one_state_loop = 1'b0;
    assign seq_loop_intf_125.one_state_block = 1'b0;
    assign seq_loop_intf_125.finish = finish;
    csv_file_dump seq_loop_csv_dumper_125;
    seq_loop_monitor #(452) seq_loop_monitor_125;
    seq_loop_intf#(452) seq_loop_intf_126(clock,reset);
    assign seq_loop_intf_126.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state395;
    assign seq_loop_intf_126.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_126.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_126.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_126.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state403;
    assign seq_loop_intf_126.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_126.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state452;
    assign seq_loop_intf_126.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_126.post_loop_state2 = 452'h0;
    assign seq_loop_intf_126.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_126.post_loop_state3 = 452'h0;
    assign seq_loop_intf_126.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_126.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state398;
    assign seq_loop_intf_126.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_126.quit_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state400;
    assign seq_loop_intf_126.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_126.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_126.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state398;
    assign seq_loop_intf_126.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state402;
    assign seq_loop_intf_126.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_126.iter_end_state1 = 452'h0;
    assign seq_loop_intf_126.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_126.one_state_loop = 1'b0;
    assign seq_loop_intf_126.one_state_block = 1'b0;
    assign seq_loop_intf_126.finish = finish;
    csv_file_dump seq_loop_csv_dumper_126;
    seq_loop_monitor #(452) seq_loop_monitor_126;
    seq_loop_intf#(452) seq_loop_intf_127(clock,reset);
    assign seq_loop_intf_127.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state368;
    assign seq_loop_intf_127.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_127.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_127.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_127.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state452;
    assign seq_loop_intf_127.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_127.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state443;
    assign seq_loop_intf_127.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_127.post_loop_state2 = 452'h0;
    assign seq_loop_intf_127.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_127.post_loop_state3 = 452'h0;
    assign seq_loop_intf_127.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_127.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state400;
    assign seq_loop_intf_127.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_127.quit_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state440;
    assign seq_loop_intf_127.quit_states_valid[1] = 1'b1;
    assign seq_loop_intf_127.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_127.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state370;
    assign seq_loop_intf_127.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state440;
    assign seq_loop_intf_127.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_127.iter_end_state1 = 452'h0;
    assign seq_loop_intf_127.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_127.one_state_loop = 1'b0;
    assign seq_loop_intf_127.one_state_block = 1'b0;
    assign seq_loop_intf_127.finish = finish;
    csv_file_dump seq_loop_csv_dumper_127;
    seq_loop_monitor #(452) seq_loop_monitor_127;
    seq_loop_intf#(452) seq_loop_intf_128(clock,reset);
    assign seq_loop_intf_128.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state444;
    assign seq_loop_intf_128.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_128.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_128.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_128.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state446;
    assign seq_loop_intf_128.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_128.post_loop_state1 = 452'h0;
    assign seq_loop_intf_128.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_128.post_loop_state2 = 452'h0;
    assign seq_loop_intf_128.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_128.post_loop_state3 = 452'h0;
    assign seq_loop_intf_128.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_128.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state445;
    assign seq_loop_intf_128.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_128.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_128.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_128.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_128.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state445;
    assign seq_loop_intf_128.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state445;
    assign seq_loop_intf_128.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_128.iter_end_state1 = 452'h0;
    assign seq_loop_intf_128.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_128.one_state_loop = 1'b1;
    assign seq_loop_intf_128.one_state_block = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state445_blk;
    assign seq_loop_intf_128.finish = finish;
    csv_file_dump seq_loop_csv_dumper_128;
    seq_loop_monitor #(452) seq_loop_monitor_128;
    seq_loop_intf#(452) seq_loop_intf_129(clock,reset);
    assign seq_loop_intf_129.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state446;
    assign seq_loop_intf_129.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_129.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_129.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_129.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state443;
    assign seq_loop_intf_129.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_129.post_loop_state1 = 452'h0;
    assign seq_loop_intf_129.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_129.post_loop_state2 = 452'h0;
    assign seq_loop_intf_129.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_129.post_loop_state3 = 452'h0;
    assign seq_loop_intf_129.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_129.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state447;
    assign seq_loop_intf_129.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_129.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_129.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_129.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_129.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state447;
    assign seq_loop_intf_129.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state447;
    assign seq_loop_intf_129.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_129.iter_end_state1 = 452'h0;
    assign seq_loop_intf_129.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_129.one_state_loop = 1'b1;
    assign seq_loop_intf_129.one_state_block = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state447_blk;
    assign seq_loop_intf_129.finish = finish;
    csv_file_dump seq_loop_csv_dumper_129;
    seq_loop_monitor #(452) seq_loop_monitor_129;
    seq_loop_intf#(452) seq_loop_intf_130(clock,reset);
    assign seq_loop_intf_130.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state440;
    assign seq_loop_intf_130.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_130.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_130.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_130.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state448;
    assign seq_loop_intf_130.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_130.post_loop_state1 = 452'h0;
    assign seq_loop_intf_130.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_130.post_loop_state2 = 452'h0;
    assign seq_loop_intf_130.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_130.post_loop_state3 = 452'h0;
    assign seq_loop_intf_130.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_130.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state443;
    assign seq_loop_intf_130.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_130.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_130.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_130.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_130.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state443;
    assign seq_loop_intf_130.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state447;
    assign seq_loop_intf_130.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_130.iter_end_state1 = 452'h0;
    assign seq_loop_intf_130.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_130.one_state_loop = 1'b0;
    assign seq_loop_intf_130.one_state_block = 1'b0;
    assign seq_loop_intf_130.finish = finish;
    csv_file_dump seq_loop_csv_dumper_130;
    seq_loop_monitor #(452) seq_loop_monitor_130;
    seq_loop_intf#(452) seq_loop_intf_131(clock,reset);
    assign seq_loop_intf_131.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state449;
    assign seq_loop_intf_131.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_131.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_131.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_131.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state449;
    assign seq_loop_intf_131.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_131.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state448;
    assign seq_loop_intf_131.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_131.post_loop_state2 = 452'h0;
    assign seq_loop_intf_131.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_131.post_loop_state3 = 452'h0;
    assign seq_loop_intf_131.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_131.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state450;
    assign seq_loop_intf_131.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_131.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_131.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_131.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_131.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state450;
    assign seq_loop_intf_131.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state451;
    assign seq_loop_intf_131.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_131.iter_end_state1 = 452'h0;
    assign seq_loop_intf_131.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_131.one_state_loop = 1'b0;
    assign seq_loop_intf_131.one_state_block = 1'b0;
    assign seq_loop_intf_131.finish = finish;
    csv_file_dump seq_loop_csv_dumper_131;
    seq_loop_monitor #(452) seq_loop_monitor_131;
    seq_loop_intf#(452) seq_loop_intf_132(clock,reset);
    assign seq_loop_intf_132.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state448;
    assign seq_loop_intf_132.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_132.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_132.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_132.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state451;
    assign seq_loop_intf_132.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_132.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state448;
    assign seq_loop_intf_132.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_132.post_loop_state2 = 452'h0;
    assign seq_loop_intf_132.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_132.post_loop_state3 = 452'h0;
    assign seq_loop_intf_132.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_132.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state450;
    assign seq_loop_intf_132.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_132.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_132.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_132.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_132.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state449;
    assign seq_loop_intf_132.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state450;
    assign seq_loop_intf_132.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_132.iter_end_state1 = 452'h0;
    assign seq_loop_intf_132.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_132.one_state_loop = 1'b0;
    assign seq_loop_intf_132.one_state_block = 1'b0;
    assign seq_loop_intf_132.finish = finish;
    csv_file_dump seq_loop_csv_dumper_132;
    seq_loop_monitor #(452) seq_loop_monitor_132;
    seq_loop_intf#(452) seq_loop_intf_133(clock,reset);
    assign seq_loop_intf_133.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state443;
    assign seq_loop_intf_133.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_133.pre_loop_state1 = 452'h0;
    assign seq_loop_intf_133.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_133.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state452;
    assign seq_loop_intf_133.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_133.post_loop_state1 = 452'h0;
    assign seq_loop_intf_133.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_133.post_loop_state2 = 452'h0;
    assign seq_loop_intf_133.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_133.post_loop_state3 = 452'h0;
    assign seq_loop_intf_133.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_133.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state448;
    assign seq_loop_intf_133.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_133.quit_loop_state1 = 452'h0;
    assign seq_loop_intf_133.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_133.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_CS_fsm;
    assign seq_loop_intf_133.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state448;
    assign seq_loop_intf_133.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.ap_ST_fsm_state450;
    assign seq_loop_intf_133.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_133.iter_end_state1 = 452'h0;
    assign seq_loop_intf_133.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_133.one_state_loop = 1'b0;
    assign seq_loop_intf_133.one_state_block = 1'b0;
    assign seq_loop_intf_133.finish = finish;
    csv_file_dump seq_loop_csv_dumper_133;
    seq_loop_monitor #(452) seq_loop_monitor_133;
    seq_loop_intf#(10) seq_loop_intf_134(clock,reset);
    assign seq_loop_intf_134.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state4;
    assign seq_loop_intf_134.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_134.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_134.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_134.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state6;
    assign seq_loop_intf_134.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_134.post_loop_state1 = 10'h0;
    assign seq_loop_intf_134.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_134.post_loop_state2 = 10'h0;
    assign seq_loop_intf_134.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_134.post_loop_state3 = 10'h0;
    assign seq_loop_intf_134.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_134.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state5;
    assign seq_loop_intf_134.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_134.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_134.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_134.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_CS_fsm;
    assign seq_loop_intf_134.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state5;
    assign seq_loop_intf_134.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state5;
    assign seq_loop_intf_134.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_134.iter_end_state1 = 10'h0;
    assign seq_loop_intf_134.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_134.one_state_loop = 1'b1;
    assign seq_loop_intf_134.one_state_block = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state5_blk;
    assign seq_loop_intf_134.finish = finish;
    csv_file_dump seq_loop_csv_dumper_134;
    seq_loop_monitor #(10) seq_loop_monitor_134;
    seq_loop_intf#(10) seq_loop_intf_135(clock,reset);
    assign seq_loop_intf_135.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state5;
    assign seq_loop_intf_135.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_135.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_135.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_135.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state8;
    assign seq_loop_intf_135.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_135.post_loop_state1 = 10'h0;
    assign seq_loop_intf_135.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_135.post_loop_state2 = 10'h0;
    assign seq_loop_intf_135.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_135.post_loop_state3 = 10'h0;
    assign seq_loop_intf_135.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_135.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state6;
    assign seq_loop_intf_135.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_135.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_135.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_135.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_CS_fsm;
    assign seq_loop_intf_135.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state6;
    assign seq_loop_intf_135.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state7;
    assign seq_loop_intf_135.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_135.iter_end_state1 = 10'h0;
    assign seq_loop_intf_135.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_135.one_state_loop = 1'b0;
    assign seq_loop_intf_135.one_state_block = 1'b0;
    assign seq_loop_intf_135.finish = finish;
    csv_file_dump seq_loop_csv_dumper_135;
    seq_loop_monitor #(10) seq_loop_monitor_135;
    seq_loop_intf#(10) seq_loop_intf_136(clock,reset);
    assign seq_loop_intf_136.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state6;
    assign seq_loop_intf_136.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_136.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_136.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_136.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state1;
    assign seq_loop_intf_136.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_136.post_loop_state1 = 10'h0;
    assign seq_loop_intf_136.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_136.post_loop_state2 = 10'h0;
    assign seq_loop_intf_136.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_136.post_loop_state3 = 10'h0;
    assign seq_loop_intf_136.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_136.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state8;
    assign seq_loop_intf_136.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_136.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_136.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_136.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_CS_fsm;
    assign seq_loop_intf_136.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state8;
    assign seq_loop_intf_136.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_mkgm2_1_fu_3306.ap_ST_fsm_state10;
    assign seq_loop_intf_136.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_136.iter_end_state1 = 10'h0;
    assign seq_loop_intf_136.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_136.one_state_loop = 1'b0;
    assign seq_loop_intf_136.one_state_block = 1'b0;
    assign seq_loop_intf_136.finish = finish;
    csv_file_dump seq_loop_csv_dumper_136;
    seq_loop_monitor #(10) seq_loop_monitor_136;
    seq_loop_intf#(14) seq_loop_intf_137(clock,reset);
    assign seq_loop_intf_137.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state1;
    assign seq_loop_intf_137.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_137.pre_loop_state1 = 14'h0;
    assign seq_loop_intf_137.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_137.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state5;
    assign seq_loop_intf_137.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_137.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state7;
    assign seq_loop_intf_137.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_137.post_loop_state2 = 14'h0;
    assign seq_loop_intf_137.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_137.post_loop_state3 = 14'h0;
    assign seq_loop_intf_137.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_137.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state2;
    assign seq_loop_intf_137.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_137.quit_loop_state1 = 14'h0;
    assign seq_loop_intf_137.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_137.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_CS_fsm;
    assign seq_loop_intf_137.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state2;
    assign seq_loop_intf_137.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state4;
    assign seq_loop_intf_137.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_137.iter_end_state1 = 14'h0;
    assign seq_loop_intf_137.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_137.one_state_loop = 1'b0;
    assign seq_loop_intf_137.one_state_block = 1'b0;
    assign seq_loop_intf_137.finish = finish;
    csv_file_dump seq_loop_csv_dumper_137;
    seq_loop_monitor #(14) seq_loop_monitor_137;
    seq_loop_intf#(14) seq_loop_intf_138(clock,reset);
    assign seq_loop_intf_138.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state2;
    assign seq_loop_intf_138.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_138.pre_loop_state1 = 14'h0;
    assign seq_loop_intf_138.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_138.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state9;
    assign seq_loop_intf_138.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_138.post_loop_state1 = 14'h0;
    assign seq_loop_intf_138.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_138.post_loop_state2 = 14'h0;
    assign seq_loop_intf_138.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_138.post_loop_state3 = 14'h0;
    assign seq_loop_intf_138.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_138.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state7;
    assign seq_loop_intf_138.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_138.quit_loop_state1 = 14'h0;
    assign seq_loop_intf_138.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_138.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_CS_fsm;
    assign seq_loop_intf_138.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state7;
    assign seq_loop_intf_138.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state8;
    assign seq_loop_intf_138.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_138.iter_end_state1 = 14'h0;
    assign seq_loop_intf_138.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_138.one_state_loop = 1'b0;
    assign seq_loop_intf_138.one_state_block = 1'b0;
    assign seq_loop_intf_138.finish = finish;
    csv_file_dump seq_loop_csv_dumper_138;
    seq_loop_monitor #(14) seq_loop_monitor_138;
    seq_loop_intf#(14) seq_loop_intf_139(clock,reset);
    assign seq_loop_intf_139.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state7;
    assign seq_loop_intf_139.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_139.pre_loop_state1 = 14'h0;
    assign seq_loop_intf_139.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_139.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state12;
    assign seq_loop_intf_139.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_139.post_loop_state1 = 14'h0;
    assign seq_loop_intf_139.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_139.post_loop_state2 = 14'h0;
    assign seq_loop_intf_139.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_139.post_loop_state3 = 14'h0;
    assign seq_loop_intf_139.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_139.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state9;
    assign seq_loop_intf_139.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_139.quit_loop_state1 = 14'h0;
    assign seq_loop_intf_139.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_139.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_CS_fsm;
    assign seq_loop_intf_139.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state9;
    assign seq_loop_intf_139.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state11;
    assign seq_loop_intf_139.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_139.iter_end_state1 = 14'h0;
    assign seq_loop_intf_139.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_139.one_state_loop = 1'b0;
    assign seq_loop_intf_139.one_state_block = 1'b0;
    assign seq_loop_intf_139.finish = finish;
    csv_file_dump seq_loop_csv_dumper_139;
    seq_loop_monitor #(14) seq_loop_monitor_139;
    seq_loop_intf#(14) seq_loop_intf_140(clock,reset);
    assign seq_loop_intf_140.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state2;
    assign seq_loop_intf_140.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_140.pre_loop_state1 = 14'h0;
    assign seq_loop_intf_140.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_140.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state14;
    assign seq_loop_intf_140.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_140.post_loop_state1 = 14'h0;
    assign seq_loop_intf_140.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_140.post_loop_state2 = 14'h0;
    assign seq_loop_intf_140.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_140.post_loop_state3 = 14'h0;
    assign seq_loop_intf_140.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_140.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state5;
    assign seq_loop_intf_140.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_140.quit_loop_state1 = 14'h0;
    assign seq_loop_intf_140.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_140.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_CS_fsm;
    assign seq_loop_intf_140.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state5;
    assign seq_loop_intf_140.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.ap_ST_fsm_state6;
    assign seq_loop_intf_140.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_140.iter_end_state1 = 14'h0;
    assign seq_loop_intf_140.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_140.one_state_loop = 1'b0;
    assign seq_loop_intf_140.one_state_block = 1'b0;
    assign seq_loop_intf_140.finish = finish;
    csv_file_dump seq_loop_csv_dumper_140;
    seq_loop_monitor #(14) seq_loop_monitor_140;
    seq_loop_intf#(60) seq_loop_intf_141(clock,reset);
    assign seq_loop_intf_141.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state2;
    assign seq_loop_intf_141.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_141.pre_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state3;
    assign seq_loop_intf_141.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_141.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state3;
    assign seq_loop_intf_141.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_141.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state6;
    assign seq_loop_intf_141.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_141.post_loop_state2 = 60'h0;
    assign seq_loop_intf_141.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_141.post_loop_state3 = 60'h0;
    assign seq_loop_intf_141.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_141.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state4;
    assign seq_loop_intf_141.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_141.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_141.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_141.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_141.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state4;
    assign seq_loop_intf_141.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state5;
    assign seq_loop_intf_141.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_141.iter_end_state1 = 60'h0;
    assign seq_loop_intf_141.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_141.one_state_loop = 1'b0;
    assign seq_loop_intf_141.one_state_block = 1'b0;
    assign seq_loop_intf_141.finish = finish;
    csv_file_dump seq_loop_csv_dumper_141;
    seq_loop_monitor #(60) seq_loop_monitor_141;
    seq_loop_intf#(60) seq_loop_intf_142(clock,reset);
    assign seq_loop_intf_142.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state2;
    assign seq_loop_intf_142.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_142.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_142.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_142.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state5;
    assign seq_loop_intf_142.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_142.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state6;
    assign seq_loop_intf_142.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_142.post_loop_state2 = 60'h0;
    assign seq_loop_intf_142.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_142.post_loop_state3 = 60'h0;
    assign seq_loop_intf_142.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_142.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state4;
    assign seq_loop_intf_142.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_142.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_142.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_142.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_142.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state3;
    assign seq_loop_intf_142.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state4;
    assign seq_loop_intf_142.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_142.iter_end_state1 = 60'h0;
    assign seq_loop_intf_142.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_142.one_state_loop = 1'b0;
    assign seq_loop_intf_142.one_state_block = 1'b0;
    assign seq_loop_intf_142.finish = finish;
    csv_file_dump seq_loop_csv_dumper_142;
    seq_loop_monitor #(60) seq_loop_monitor_142;
    seq_loop_intf#(60) seq_loop_intf_143(clock,reset);
    assign seq_loop_intf_143.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state10;
    assign seq_loop_intf_143.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_143.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_143.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_143.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state13;
    assign seq_loop_intf_143.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_143.post_loop_state1 = 60'h0;
    assign seq_loop_intf_143.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_143.post_loop_state2 = 60'h0;
    assign seq_loop_intf_143.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_143.post_loop_state3 = 60'h0;
    assign seq_loop_intf_143.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_143.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state11;
    assign seq_loop_intf_143.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_143.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_143.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_143.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_143.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state11;
    assign seq_loop_intf_143.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state12;
    assign seq_loop_intf_143.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_143.iter_end_state1 = 60'h0;
    assign seq_loop_intf_143.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_143.one_state_loop = 1'b0;
    assign seq_loop_intf_143.one_state_block = 1'b0;
    assign seq_loop_intf_143.finish = finish;
    csv_file_dump seq_loop_csv_dumper_143;
    seq_loop_monitor #(60) seq_loop_monitor_143;
    seq_loop_intf#(60) seq_loop_intf_144(clock,reset);
    assign seq_loop_intf_144.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state14;
    assign seq_loop_intf_144.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_144.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_144.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_144.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state18;
    assign seq_loop_intf_144.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_144.post_loop_state1 = 60'h0;
    assign seq_loop_intf_144.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_144.post_loop_state2 = 60'h0;
    assign seq_loop_intf_144.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_144.post_loop_state3 = 60'h0;
    assign seq_loop_intf_144.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_144.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state15;
    assign seq_loop_intf_144.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_144.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_144.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_144.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_144.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state15;
    assign seq_loop_intf_144.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state17;
    assign seq_loop_intf_144.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_144.iter_end_state1 = 60'h0;
    assign seq_loop_intf_144.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_144.one_state_loop = 1'b0;
    assign seq_loop_intf_144.one_state_block = 1'b0;
    assign seq_loop_intf_144.finish = finish;
    csv_file_dump seq_loop_csv_dumper_144;
    seq_loop_monitor #(60) seq_loop_monitor_144;
    seq_loop_intf#(60) seq_loop_intf_145(clock,reset);
    assign seq_loop_intf_145.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state18;
    assign seq_loop_intf_145.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_145.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_145.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_145.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state21;
    assign seq_loop_intf_145.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_145.post_loop_state1 = 60'h0;
    assign seq_loop_intf_145.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_145.post_loop_state2 = 60'h0;
    assign seq_loop_intf_145.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_145.post_loop_state3 = 60'h0;
    assign seq_loop_intf_145.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_145.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state19;
    assign seq_loop_intf_145.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_145.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_145.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_145.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_145.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state19;
    assign seq_loop_intf_145.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state20;
    assign seq_loop_intf_145.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_145.iter_end_state1 = 60'h0;
    assign seq_loop_intf_145.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_145.one_state_loop = 1'b0;
    assign seq_loop_intf_145.one_state_block = 1'b0;
    assign seq_loop_intf_145.finish = finish;
    csv_file_dump seq_loop_csv_dumper_145;
    seq_loop_monitor #(60) seq_loop_monitor_145;
    seq_loop_intf#(60) seq_loop_intf_146(clock,reset);
    assign seq_loop_intf_146.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state21;
    assign seq_loop_intf_146.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_146.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_146.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_146.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state25;
    assign seq_loop_intf_146.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_146.post_loop_state1 = 60'h0;
    assign seq_loop_intf_146.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_146.post_loop_state2 = 60'h0;
    assign seq_loop_intf_146.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_146.post_loop_state3 = 60'h0;
    assign seq_loop_intf_146.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_146.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state22;
    assign seq_loop_intf_146.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_146.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_146.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_146.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_146.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state22;
    assign seq_loop_intf_146.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state24;
    assign seq_loop_intf_146.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_146.iter_end_state1 = 60'h0;
    assign seq_loop_intf_146.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_146.one_state_loop = 1'b0;
    assign seq_loop_intf_146.one_state_block = 1'b0;
    assign seq_loop_intf_146.finish = finish;
    csv_file_dump seq_loop_csv_dumper_146;
    seq_loop_monitor #(60) seq_loop_monitor_146;
    seq_loop_intf#(60) seq_loop_intf_147(clock,reset);
    assign seq_loop_intf_147.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state4;
    assign seq_loop_intf_147.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_147.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_147.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_147.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state30;
    assign seq_loop_intf_147.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_147.post_loop_state1 = 60'h0;
    assign seq_loop_intf_147.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_147.post_loop_state2 = 60'h0;
    assign seq_loop_intf_147.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_147.post_loop_state3 = 60'h0;
    assign seq_loop_intf_147.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_147.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state6;
    assign seq_loop_intf_147.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_147.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_147.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_147.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_147.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state6;
    assign seq_loop_intf_147.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state29;
    assign seq_loop_intf_147.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_147.iter_end_state1 = 60'h0;
    assign seq_loop_intf_147.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_147.one_state_loop = 1'b0;
    assign seq_loop_intf_147.one_state_block = 1'b0;
    assign seq_loop_intf_147.finish = finish;
    csv_file_dump seq_loop_csv_dumper_147;
    seq_loop_monitor #(60) seq_loop_monitor_147;
    seq_loop_intf#(60) seq_loop_intf_148(clock,reset);
    assign seq_loop_intf_148.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state37;
    assign seq_loop_intf_148.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_148.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_148.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_148.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state40;
    assign seq_loop_intf_148.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_148.post_loop_state1 = 60'h0;
    assign seq_loop_intf_148.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_148.post_loop_state2 = 60'h0;
    assign seq_loop_intf_148.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_148.post_loop_state3 = 60'h0;
    assign seq_loop_intf_148.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_148.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state38;
    assign seq_loop_intf_148.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_148.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_148.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_148.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_148.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state38;
    assign seq_loop_intf_148.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state39;
    assign seq_loop_intf_148.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_148.iter_end_state1 = 60'h0;
    assign seq_loop_intf_148.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_148.one_state_loop = 1'b0;
    assign seq_loop_intf_148.one_state_block = 1'b0;
    assign seq_loop_intf_148.finish = finish;
    csv_file_dump seq_loop_csv_dumper_148;
    seq_loop_monitor #(60) seq_loop_monitor_148;
    seq_loop_intf#(60) seq_loop_intf_149(clock,reset);
    assign seq_loop_intf_149.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state42;
    assign seq_loop_intf_149.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_149.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_149.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_149.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state45;
    assign seq_loop_intf_149.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_149.post_loop_state1 = 60'h0;
    assign seq_loop_intf_149.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_149.post_loop_state2 = 60'h0;
    assign seq_loop_intf_149.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_149.post_loop_state3 = 60'h0;
    assign seq_loop_intf_149.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_149.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state44;
    assign seq_loop_intf_149.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_149.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_149.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_149.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_149.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state43;
    assign seq_loop_intf_149.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state44;
    assign seq_loop_intf_149.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_149.iter_end_state1 = 60'h0;
    assign seq_loop_intf_149.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_149.one_state_loop = 1'b0;
    assign seq_loop_intf_149.one_state_block = 1'b0;
    assign seq_loop_intf_149.finish = finish;
    csv_file_dump seq_loop_csv_dumper_149;
    seq_loop_monitor #(60) seq_loop_monitor_149;
    seq_loop_intf#(60) seq_loop_intf_150(clock,reset);
    assign seq_loop_intf_150.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state41;
    assign seq_loop_intf_150.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_150.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_150.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_150.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state46;
    assign seq_loop_intf_150.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_150.post_loop_state1 = 60'h0;
    assign seq_loop_intf_150.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_150.post_loop_state2 = 60'h0;
    assign seq_loop_intf_150.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_150.post_loop_state3 = 60'h0;
    assign seq_loop_intf_150.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_150.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state42;
    assign seq_loop_intf_150.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_150.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_150.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_150.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_150.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state42;
    assign seq_loop_intf_150.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state45;
    assign seq_loop_intf_150.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_150.iter_end_state1 = 60'h0;
    assign seq_loop_intf_150.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_150.one_state_loop = 1'b0;
    assign seq_loop_intf_150.one_state_block = 1'b0;
    assign seq_loop_intf_150.finish = finish;
    csv_file_dump seq_loop_csv_dumper_150;
    seq_loop_monitor #(60) seq_loop_monitor_150;
    seq_loop_intf#(60) seq_loop_intf_151(clock,reset);
    assign seq_loop_intf_151.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state46;
    assign seq_loop_intf_151.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_151.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_151.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_151.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state50;
    assign seq_loop_intf_151.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_151.post_loop_state1 = 60'h0;
    assign seq_loop_intf_151.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_151.post_loop_state2 = 60'h0;
    assign seq_loop_intf_151.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_151.post_loop_state3 = 60'h0;
    assign seq_loop_intf_151.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_151.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state47;
    assign seq_loop_intf_151.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_151.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_151.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_151.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_151.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state47;
    assign seq_loop_intf_151.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state49;
    assign seq_loop_intf_151.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_151.iter_end_state1 = 60'h0;
    assign seq_loop_intf_151.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_151.one_state_loop = 1'b0;
    assign seq_loop_intf_151.one_state_block = 1'b0;
    assign seq_loop_intf_151.finish = finish;
    csv_file_dump seq_loop_csv_dumper_151;
    seq_loop_monitor #(60) seq_loop_monitor_151;
    seq_loop_intf#(60) seq_loop_intf_152(clock,reset);
    assign seq_loop_intf_152.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state50;
    assign seq_loop_intf_152.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_152.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_152.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_152.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state53;
    assign seq_loop_intf_152.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_152.post_loop_state1 = 60'h0;
    assign seq_loop_intf_152.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_152.post_loop_state2 = 60'h0;
    assign seq_loop_intf_152.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_152.post_loop_state3 = 60'h0;
    assign seq_loop_intf_152.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_152.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state52;
    assign seq_loop_intf_152.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_152.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_152.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_152.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_152.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state51;
    assign seq_loop_intf_152.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state52;
    assign seq_loop_intf_152.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_152.iter_end_state1 = 60'h0;
    assign seq_loop_intf_152.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_152.one_state_loop = 1'b0;
    assign seq_loop_intf_152.one_state_block = 1'b0;
    assign seq_loop_intf_152.finish = finish;
    csv_file_dump seq_loop_csv_dumper_152;
    seq_loop_monitor #(60) seq_loop_monitor_152;
    seq_loop_intf#(60) seq_loop_intf_153(clock,reset);
    assign seq_loop_intf_153.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state47;
    assign seq_loop_intf_153.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_153.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_153.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_153.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state54;
    assign seq_loop_intf_153.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_153.post_loop_state1 = 60'h0;
    assign seq_loop_intf_153.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_153.post_loop_state2 = 60'h0;
    assign seq_loop_intf_153.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_153.post_loop_state3 = 60'h0;
    assign seq_loop_intf_153.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_153.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state50;
    assign seq_loop_intf_153.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_153.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_153.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_153.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_153.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state50;
    assign seq_loop_intf_153.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state53;
    assign seq_loop_intf_153.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_153.iter_end_state1 = 60'h0;
    assign seq_loop_intf_153.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_153.one_state_loop = 1'b0;
    assign seq_loop_intf_153.one_state_block = 1'b0;
    assign seq_loop_intf_153.finish = finish;
    csv_file_dump seq_loop_csv_dumper_153;
    seq_loop_monitor #(60) seq_loop_monitor_153;
    seq_loop_intf#(60) seq_loop_intf_154(clock,reset);
    assign seq_loop_intf_154.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state54;
    assign seq_loop_intf_154.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_154.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_154.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_154.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state58;
    assign seq_loop_intf_154.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_154.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state60;
    assign seq_loop_intf_154.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_154.post_loop_state2 = 60'h0;
    assign seq_loop_intf_154.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_154.post_loop_state3 = 60'h0;
    assign seq_loop_intf_154.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_154.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state55;
    assign seq_loop_intf_154.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_154.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_154.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_154.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_154.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state55;
    assign seq_loop_intf_154.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state57;
    assign seq_loop_intf_154.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_154.iter_end_state1 = 60'h0;
    assign seq_loop_intf_154.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_154.one_state_loop = 1'b0;
    assign seq_loop_intf_154.one_state_block = 1'b0;
    assign seq_loop_intf_154.finish = finish;
    csv_file_dump seq_loop_csv_dumper_154;
    seq_loop_monitor #(60) seq_loop_monitor_154;
    seq_loop_intf#(60) seq_loop_intf_155(clock,reset);
    assign seq_loop_intf_155.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state32;
    assign seq_loop_intf_155.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_155.pre_loop_state1 = 60'h0;
    assign seq_loop_intf_155.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_155.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state1;
    assign seq_loop_intf_155.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_155.post_loop_state1 = 60'h0;
    assign seq_loop_intf_155.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_155.post_loop_state2 = 60'h0;
    assign seq_loop_intf_155.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_155.post_loop_state3 = 60'h0;
    assign seq_loop_intf_155.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_155.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state33;
    assign seq_loop_intf_155.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_155.quit_loop_state1 = 60'h0;
    assign seq_loop_intf_155.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_155.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_CS_fsm;
    assign seq_loop_intf_155.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state33;
    assign seq_loop_intf_155.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.ap_ST_fsm_state60;
    assign seq_loop_intf_155.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_155.iter_end_state1 = 60'h0;
    assign seq_loop_intf_155.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_155.one_state_loop = 1'b0;
    assign seq_loop_intf_155.one_state_block = 1'b0;
    assign seq_loop_intf_155.finish = finish;
    csv_file_dump seq_loop_csv_dumper_155;
    seq_loop_monitor #(60) seq_loop_monitor_155;
    seq_loop_intf#(19) seq_loop_intf_156(clock,reset);
    assign seq_loop_intf_156.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state8;
    assign seq_loop_intf_156.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_156.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_156.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_156.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state11;
    assign seq_loop_intf_156.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_156.post_loop_state1 = 19'h0;
    assign seq_loop_intf_156.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_156.post_loop_state2 = 19'h0;
    assign seq_loop_intf_156.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_156.post_loop_state3 = 19'h0;
    assign seq_loop_intf_156.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_156.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state10;
    assign seq_loop_intf_156.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_156.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_156.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_156.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_CS_fsm;
    assign seq_loop_intf_156.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state9;
    assign seq_loop_intf_156.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state10;
    assign seq_loop_intf_156.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_156.iter_end_state1 = 19'h0;
    assign seq_loop_intf_156.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_156.one_state_loop = 1'b0;
    assign seq_loop_intf_156.one_state_block = 1'b0;
    assign seq_loop_intf_156.finish = finish;
    csv_file_dump seq_loop_csv_dumper_156;
    seq_loop_monitor #(19) seq_loop_monitor_156;
    seq_loop_intf#(19) seq_loop_intf_157(clock,reset);
    assign seq_loop_intf_157.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state10;
    assign seq_loop_intf_157.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_157.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_157.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_157.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state7;
    assign seq_loop_intf_157.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_157.post_loop_state1 = 19'h0;
    assign seq_loop_intf_157.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_157.post_loop_state2 = 19'h0;
    assign seq_loop_intf_157.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_157.post_loop_state3 = 19'h0;
    assign seq_loop_intf_157.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_157.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state11;
    assign seq_loop_intf_157.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_157.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_157.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_157.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_CS_fsm;
    assign seq_loop_intf_157.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state11;
    assign seq_loop_intf_157.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state12;
    assign seq_loop_intf_157.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_157.iter_end_state1 = 19'h0;
    assign seq_loop_intf_157.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_157.one_state_loop = 1'b0;
    assign seq_loop_intf_157.one_state_block = 1'b0;
    assign seq_loop_intf_157.finish = finish;
    csv_file_dump seq_loop_csv_dumper_157;
    seq_loop_monitor #(19) seq_loop_monitor_157;
    seq_loop_intf#(19) seq_loop_intf_158(clock,reset);
    assign seq_loop_intf_158.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state6;
    assign seq_loop_intf_158.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_158.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_158.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_158.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state13;
    assign seq_loop_intf_158.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_158.post_loop_state1 = 19'h0;
    assign seq_loop_intf_158.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_158.post_loop_state2 = 19'h0;
    assign seq_loop_intf_158.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_158.post_loop_state3 = 19'h0;
    assign seq_loop_intf_158.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_158.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state7;
    assign seq_loop_intf_158.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_158.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_158.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_158.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_CS_fsm;
    assign seq_loop_intf_158.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state7;
    assign seq_loop_intf_158.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state11;
    assign seq_loop_intf_158.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_158.iter_end_state1 = 19'h0;
    assign seq_loop_intf_158.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_158.one_state_loop = 1'b0;
    assign seq_loop_intf_158.one_state_block = 1'b0;
    assign seq_loop_intf_158.finish = finish;
    csv_file_dump seq_loop_csv_dumper_158;
    seq_loop_monitor #(19) seq_loop_monitor_158;
    seq_loop_intf#(19) seq_loop_intf_159(clock,reset);
    assign seq_loop_intf_159.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state7;
    assign seq_loop_intf_159.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_159.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_159.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_159.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state2;
    assign seq_loop_intf_159.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_159.post_loop_state1 = 19'h0;
    assign seq_loop_intf_159.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_159.post_loop_state2 = 19'h0;
    assign seq_loop_intf_159.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_159.post_loop_state3 = 19'h0;
    assign seq_loop_intf_159.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_159.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state13;
    assign seq_loop_intf_159.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_159.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_159.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_159.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_CS_fsm;
    assign seq_loop_intf_159.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state13;
    assign seq_loop_intf_159.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state14;
    assign seq_loop_intf_159.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_159.iter_end_state1 = 19'h0;
    assign seq_loop_intf_159.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_159.one_state_loop = 1'b0;
    assign seq_loop_intf_159.one_state_block = 1'b0;
    assign seq_loop_intf_159.finish = finish;
    csv_file_dump seq_loop_csv_dumper_159;
    seq_loop_monitor #(19) seq_loop_monitor_159;
    seq_loop_intf#(19) seq_loop_intf_160(clock,reset);
    assign seq_loop_intf_160.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state1;
    assign seq_loop_intf_160.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_160.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_160.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_160.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state15;
    assign seq_loop_intf_160.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_160.post_loop_state1 = 19'h0;
    assign seq_loop_intf_160.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_160.post_loop_state2 = 19'h0;
    assign seq_loop_intf_160.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_160.post_loop_state3 = 19'h0;
    assign seq_loop_intf_160.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_160.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state2;
    assign seq_loop_intf_160.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_160.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_160.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_160.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_CS_fsm;
    assign seq_loop_intf_160.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state2;
    assign seq_loop_intf_160.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state13;
    assign seq_loop_intf_160.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_160.iter_end_state1 = 19'h0;
    assign seq_loop_intf_160.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_160.one_state_loop = 1'b0;
    assign seq_loop_intf_160.one_state_block = 1'b0;
    assign seq_loop_intf_160.finish = finish;
    csv_file_dump seq_loop_csv_dumper_160;
    seq_loop_monitor #(19) seq_loop_monitor_160;
    seq_loop_intf#(19) seq_loop_intf_161(clock,reset);
    assign seq_loop_intf_161.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state15;
    assign seq_loop_intf_161.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_161.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_161.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_161.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state18;
    assign seq_loop_intf_161.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_161.post_loop_state1 = 19'h0;
    assign seq_loop_intf_161.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_161.post_loop_state2 = 19'h0;
    assign seq_loop_intf_161.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_161.post_loop_state3 = 19'h0;
    assign seq_loop_intf_161.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_161.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state17;
    assign seq_loop_intf_161.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_161.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_161.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_161.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_CS_fsm;
    assign seq_loop_intf_161.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state16;
    assign seq_loop_intf_161.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state17;
    assign seq_loop_intf_161.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_161.iter_end_state1 = 19'h0;
    assign seq_loop_intf_161.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_161.one_state_loop = 1'b0;
    assign seq_loop_intf_161.one_state_block = 1'b0;
    assign seq_loop_intf_161.finish = finish;
    csv_file_dump seq_loop_csv_dumper_161;
    seq_loop_monitor #(19) seq_loop_monitor_161;
    seq_loop_intf#(19) seq_loop_intf_162(clock,reset);
    assign seq_loop_intf_162.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state17;
    assign seq_loop_intf_162.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_162.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_162.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_162.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state15;
    assign seq_loop_intf_162.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_162.post_loop_state1 = 19'h0;
    assign seq_loop_intf_162.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_162.post_loop_state2 = 19'h0;
    assign seq_loop_intf_162.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_162.post_loop_state3 = 19'h0;
    assign seq_loop_intf_162.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_162.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state18;
    assign seq_loop_intf_162.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_162.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_162.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_162.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_CS_fsm;
    assign seq_loop_intf_162.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state18;
    assign seq_loop_intf_162.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state19;
    assign seq_loop_intf_162.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_162.iter_end_state1 = 19'h0;
    assign seq_loop_intf_162.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_162.one_state_loop = 1'b0;
    assign seq_loop_intf_162.one_state_block = 1'b0;
    assign seq_loop_intf_162.finish = finish;
    csv_file_dump seq_loop_csv_dumper_162;
    seq_loop_monitor #(19) seq_loop_monitor_162;
    seq_loop_intf#(19) seq_loop_intf_163(clock,reset);
    assign seq_loop_intf_163.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state2;
    assign seq_loop_intf_163.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_163.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_163.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_163.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state1;
    assign seq_loop_intf_163.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_163.post_loop_state1 = 19'h0;
    assign seq_loop_intf_163.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_163.post_loop_state2 = 19'h0;
    assign seq_loop_intf_163.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_163.post_loop_state3 = 19'h0;
    assign seq_loop_intf_163.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_163.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state15;
    assign seq_loop_intf_163.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_163.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_163.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_163.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_CS_fsm;
    assign seq_loop_intf_163.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state15;
    assign seq_loop_intf_163.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_zint_rebuild_CRT_1_fu_780.ap_ST_fsm_state18;
    assign seq_loop_intf_163.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_163.iter_end_state1 = 19'h0;
    assign seq_loop_intf_163.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_163.one_state_loop = 1'b0;
    assign seq_loop_intf_163.one_state_block = 1'b0;
    assign seq_loop_intf_163.finish = finish;
    csv_file_dump seq_loop_csv_dumper_163;
    seq_loop_monitor #(19) seq_loop_monitor_163;
    seq_loop_intf#(10) seq_loop_intf_164(clock,reset);
    assign seq_loop_intf_164.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state4;
    assign seq_loop_intf_164.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_164.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_164.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_164.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state6;
    assign seq_loop_intf_164.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_164.post_loop_state1 = 10'h0;
    assign seq_loop_intf_164.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_164.post_loop_state2 = 10'h0;
    assign seq_loop_intf_164.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_164.post_loop_state3 = 10'h0;
    assign seq_loop_intf_164.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_164.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state5;
    assign seq_loop_intf_164.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_164.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_164.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_164.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_CS_fsm;
    assign seq_loop_intf_164.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state5;
    assign seq_loop_intf_164.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state5;
    assign seq_loop_intf_164.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_164.iter_end_state1 = 10'h0;
    assign seq_loop_intf_164.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_164.one_state_loop = 1'b1;
    assign seq_loop_intf_164.one_state_block = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state5_blk;
    assign seq_loop_intf_164.finish = finish;
    csv_file_dump seq_loop_csv_dumper_164;
    seq_loop_monitor #(10) seq_loop_monitor_164;
    seq_loop_intf#(10) seq_loop_intf_165(clock,reset);
    assign seq_loop_intf_165.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state5;
    assign seq_loop_intf_165.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_165.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_165.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_165.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state8;
    assign seq_loop_intf_165.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_165.post_loop_state1 = 10'h0;
    assign seq_loop_intf_165.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_165.post_loop_state2 = 10'h0;
    assign seq_loop_intf_165.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_165.post_loop_state3 = 10'h0;
    assign seq_loop_intf_165.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_165.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state6;
    assign seq_loop_intf_165.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_165.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_165.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_165.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_CS_fsm;
    assign seq_loop_intf_165.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state6;
    assign seq_loop_intf_165.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state7;
    assign seq_loop_intf_165.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_165.iter_end_state1 = 10'h0;
    assign seq_loop_intf_165.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_165.one_state_loop = 1'b0;
    assign seq_loop_intf_165.one_state_block = 1'b0;
    assign seq_loop_intf_165.finish = finish;
    csv_file_dump seq_loop_csv_dumper_165;
    seq_loop_monitor #(10) seq_loop_monitor_165;
    seq_loop_intf#(10) seq_loop_intf_166(clock,reset);
    assign seq_loop_intf_166.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state6;
    assign seq_loop_intf_166.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_166.pre_loop_state1 = 10'h0;
    assign seq_loop_intf_166.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_166.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state1;
    assign seq_loop_intf_166.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_166.post_loop_state1 = 10'h0;
    assign seq_loop_intf_166.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_166.post_loop_state2 = 10'h0;
    assign seq_loop_intf_166.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_166.post_loop_state3 = 10'h0;
    assign seq_loop_intf_166.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_166.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state8;
    assign seq_loop_intf_166.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_166.quit_loop_state1 = 10'h0;
    assign seq_loop_intf_166.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_166.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_CS_fsm;
    assign seq_loop_intf_166.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state8;
    assign seq_loop_intf_166.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_mkgm2_1_fu_826.ap_ST_fsm_state10;
    assign seq_loop_intf_166.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_166.iter_end_state1 = 10'h0;
    assign seq_loop_intf_166.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_166.one_state_loop = 1'b0;
    assign seq_loop_intf_166.one_state_block = 1'b0;
    assign seq_loop_intf_166.finish = finish;
    csv_file_dump seq_loop_csv_dumper_166;
    seq_loop_monitor #(10) seq_loop_monitor_166;
    seq_loop_intf#(9) seq_loop_intf_167(clock,reset);
    assign seq_loop_intf_167.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state6;
    assign seq_loop_intf_167.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_167.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_167.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_167.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state3;
    assign seq_loop_intf_167.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_167.post_loop_state1 = 9'h0;
    assign seq_loop_intf_167.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_167.post_loop_state2 = 9'h0;
    assign seq_loop_intf_167.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_167.post_loop_state3 = 9'h0;
    assign seq_loop_intf_167.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_167.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state7;
    assign seq_loop_intf_167.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_167.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_167.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_167.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_CS_fsm;
    assign seq_loop_intf_167.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state7;
    assign seq_loop_intf_167.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state9;
    assign seq_loop_intf_167.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_167.iter_end_state1 = 9'h0;
    assign seq_loop_intf_167.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_167.one_state_loop = 1'b0;
    assign seq_loop_intf_167.one_state_block = 1'b0;
    assign seq_loop_intf_167.finish = finish;
    csv_file_dump seq_loop_csv_dumper_167;
    seq_loop_monitor #(9) seq_loop_monitor_167;
    seq_loop_intf#(9) seq_loop_intf_168(clock,reset);
    assign seq_loop_intf_168.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state2;
    assign seq_loop_intf_168.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_168.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_168.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_168.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state2;
    assign seq_loop_intf_168.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_168.post_loop_state1 = 9'h0;
    assign seq_loop_intf_168.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_168.post_loop_state2 = 9'h0;
    assign seq_loop_intf_168.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_168.post_loop_state3 = 9'h0;
    assign seq_loop_intf_168.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_168.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state3;
    assign seq_loop_intf_168.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_168.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_168.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_168.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_CS_fsm;
    assign seq_loop_intf_168.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state3;
    assign seq_loop_intf_168.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state7;
    assign seq_loop_intf_168.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_168.iter_end_state1 = 9'h0;
    assign seq_loop_intf_168.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_168.one_state_loop = 1'b0;
    assign seq_loop_intf_168.one_state_block = 1'b0;
    assign seq_loop_intf_168.finish = finish;
    csv_file_dump seq_loop_csv_dumper_168;
    seq_loop_monitor #(9) seq_loop_monitor_168;
    seq_loop_intf#(9) seq_loop_intf_169(clock,reset);
    assign seq_loop_intf_169.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state1;
    assign seq_loop_intf_169.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_169.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_169.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_169.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state1;
    assign seq_loop_intf_169.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_169.post_loop_state1 = 9'h0;
    assign seq_loop_intf_169.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_169.post_loop_state2 = 9'h0;
    assign seq_loop_intf_169.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_169.post_loop_state3 = 9'h0;
    assign seq_loop_intf_169.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_169.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state2;
    assign seq_loop_intf_169.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_169.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_169.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_169.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_CS_fsm;
    assign seq_loop_intf_169.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state2;
    assign seq_loop_intf_169.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_NTT2_ext_1_fu_841.ap_ST_fsm_state3;
    assign seq_loop_intf_169.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_169.iter_end_state1 = 9'h0;
    assign seq_loop_intf_169.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_169.one_state_loop = 1'b0;
    assign seq_loop_intf_169.one_state_block = 1'b0;
    assign seq_loop_intf_169.finish = finish;
    csv_file_dump seq_loop_csv_dumper_169;
    seq_loop_monitor #(9) seq_loop_monitor_169;
    seq_loop_intf#(11) seq_loop_intf_170(clock,reset);
    assign seq_loop_intf_170.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state6;
    assign seq_loop_intf_170.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_170.pre_loop_state1 = 11'h0;
    assign seq_loop_intf_170.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_170.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state3;
    assign seq_loop_intf_170.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_170.post_loop_state1 = 11'h0;
    assign seq_loop_intf_170.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_170.post_loop_state2 = 11'h0;
    assign seq_loop_intf_170.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_170.post_loop_state3 = 11'h0;
    assign seq_loop_intf_170.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_170.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state7;
    assign seq_loop_intf_170.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_170.quit_loop_state1 = 11'h0;
    assign seq_loop_intf_170.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_170.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_CS_fsm;
    assign seq_loop_intf_170.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state7;
    assign seq_loop_intf_170.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state9;
    assign seq_loop_intf_170.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_170.iter_end_state1 = 11'h0;
    assign seq_loop_intf_170.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_170.one_state_loop = 1'b0;
    assign seq_loop_intf_170.one_state_block = 1'b0;
    assign seq_loop_intf_170.finish = finish;
    csv_file_dump seq_loop_csv_dumper_170;
    seq_loop_monitor #(11) seq_loop_monitor_170;
    seq_loop_intf#(11) seq_loop_intf_171(clock,reset);
    assign seq_loop_intf_171.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state2;
    assign seq_loop_intf_171.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_171.pre_loop_state1 = 11'h0;
    assign seq_loop_intf_171.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_171.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state2;
    assign seq_loop_intf_171.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_171.post_loop_state1 = 11'h0;
    assign seq_loop_intf_171.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_171.post_loop_state2 = 11'h0;
    assign seq_loop_intf_171.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_171.post_loop_state3 = 11'h0;
    assign seq_loop_intf_171.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_171.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state3;
    assign seq_loop_intf_171.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_171.quit_loop_state1 = 11'h0;
    assign seq_loop_intf_171.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_171.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_CS_fsm;
    assign seq_loop_intf_171.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state3;
    assign seq_loop_intf_171.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state7;
    assign seq_loop_intf_171.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_171.iter_end_state1 = 11'h0;
    assign seq_loop_intf_171.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_171.one_state_loop = 1'b0;
    assign seq_loop_intf_171.one_state_block = 1'b0;
    assign seq_loop_intf_171.finish = finish;
    csv_file_dump seq_loop_csv_dumper_171;
    seq_loop_monitor #(11) seq_loop_monitor_171;
    seq_loop_intf#(11) seq_loop_intf_172(clock,reset);
    assign seq_loop_intf_172.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state1;
    assign seq_loop_intf_172.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_172.pre_loop_state1 = 11'h0;
    assign seq_loop_intf_172.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_172.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state10;
    assign seq_loop_intf_172.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_172.post_loop_state1 = 11'h0;
    assign seq_loop_intf_172.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_172.post_loop_state2 = 11'h0;
    assign seq_loop_intf_172.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_172.post_loop_state3 = 11'h0;
    assign seq_loop_intf_172.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_172.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state2;
    assign seq_loop_intf_172.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_172.quit_loop_state1 = 11'h0;
    assign seq_loop_intf_172.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_172.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_CS_fsm;
    assign seq_loop_intf_172.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state2;
    assign seq_loop_intf_172.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state3;
    assign seq_loop_intf_172.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_172.iter_end_state1 = 11'h0;
    assign seq_loop_intf_172.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_172.one_state_loop = 1'b0;
    assign seq_loop_intf_172.one_state_block = 1'b0;
    assign seq_loop_intf_172.finish = finish;
    csv_file_dump seq_loop_csv_dumper_172;
    seq_loop_monitor #(11) seq_loop_monitor_172;
    seq_loop_intf#(11) seq_loop_intf_173(clock,reset);
    assign seq_loop_intf_173.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state1;
    assign seq_loop_intf_173.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_173.pre_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state2;
    assign seq_loop_intf_173.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_173.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state1;
    assign seq_loop_intf_173.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_173.post_loop_state1 = 11'h0;
    assign seq_loop_intf_173.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_173.post_loop_state2 = 11'h0;
    assign seq_loop_intf_173.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_173.post_loop_state3 = 11'h0;
    assign seq_loop_intf_173.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_173.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state10;
    assign seq_loop_intf_173.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_173.quit_loop_state1 = 11'h0;
    assign seq_loop_intf_173.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_173.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_CS_fsm;
    assign seq_loop_intf_173.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state10;
    assign seq_loop_intf_173.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_make_fg_step_1_fu_234.grp_modp_iNTT2_ext_1_fu_854.ap_ST_fsm_state11;
    assign seq_loop_intf_173.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_173.iter_end_state1 = 11'h0;
    assign seq_loop_intf_173.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_173.one_state_loop = 1'b0;
    assign seq_loop_intf_173.one_state_block = 1'b0;
    assign seq_loop_intf_173.finish = finish;
    csv_file_dump seq_loop_csv_dumper_173;
    seq_loop_monitor #(11) seq_loop_monitor_173;
    seq_loop_intf#(9) seq_loop_intf_174(clock,reset);
    assign seq_loop_intf_174.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state6;
    assign seq_loop_intf_174.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_174.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_174.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_174.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state3;
    assign seq_loop_intf_174.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_174.post_loop_state1 = 9'h0;
    assign seq_loop_intf_174.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_174.post_loop_state2 = 9'h0;
    assign seq_loop_intf_174.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_174.post_loop_state3 = 9'h0;
    assign seq_loop_intf_174.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_174.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state7;
    assign seq_loop_intf_174.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_174.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_174.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_174.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_CS_fsm;
    assign seq_loop_intf_174.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state7;
    assign seq_loop_intf_174.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state9;
    assign seq_loop_intf_174.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_174.iter_end_state1 = 9'h0;
    assign seq_loop_intf_174.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_174.one_state_loop = 1'b0;
    assign seq_loop_intf_174.one_state_block = 1'b0;
    assign seq_loop_intf_174.finish = finish;
    csv_file_dump seq_loop_csv_dumper_174;
    seq_loop_monitor #(9) seq_loop_monitor_174;
    seq_loop_intf#(9) seq_loop_intf_175(clock,reset);
    assign seq_loop_intf_175.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state2;
    assign seq_loop_intf_175.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_175.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_175.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_175.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state2;
    assign seq_loop_intf_175.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_175.post_loop_state1 = 9'h0;
    assign seq_loop_intf_175.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_175.post_loop_state2 = 9'h0;
    assign seq_loop_intf_175.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_175.post_loop_state3 = 9'h0;
    assign seq_loop_intf_175.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_175.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state3;
    assign seq_loop_intf_175.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_175.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_175.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_175.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_CS_fsm;
    assign seq_loop_intf_175.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state3;
    assign seq_loop_intf_175.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state7;
    assign seq_loop_intf_175.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_175.iter_end_state1 = 9'h0;
    assign seq_loop_intf_175.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_175.one_state_loop = 1'b0;
    assign seq_loop_intf_175.one_state_block = 1'b0;
    assign seq_loop_intf_175.finish = finish;
    csv_file_dump seq_loop_csv_dumper_175;
    seq_loop_monitor #(9) seq_loop_monitor_175;
    seq_loop_intf#(9) seq_loop_intf_176(clock,reset);
    assign seq_loop_intf_176.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state1;
    assign seq_loop_intf_176.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_176.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_176.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_176.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state1;
    assign seq_loop_intf_176.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_176.post_loop_state1 = 9'h0;
    assign seq_loop_intf_176.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_176.post_loop_state2 = 9'h0;
    assign seq_loop_intf_176.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_176.post_loop_state3 = 9'h0;
    assign seq_loop_intf_176.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_176.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state2;
    assign seq_loop_intf_176.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_176.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_176.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_176.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_CS_fsm;
    assign seq_loop_intf_176.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state2;
    assign seq_loop_intf_176.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_make_fg_1_fu_3330.grp_modp_NTT2_ext_1_fu_281.ap_ST_fsm_state3;
    assign seq_loop_intf_176.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_176.iter_end_state1 = 9'h0;
    assign seq_loop_intf_176.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_176.one_state_loop = 1'b0;
    assign seq_loop_intf_176.one_state_block = 1'b0;
    assign seq_loop_intf_176.finish = finish;
    csv_file_dump seq_loop_csv_dumper_176;
    seq_loop_monitor #(9) seq_loop_monitor_176;
    seq_loop_intf#(9) seq_loop_intf_177(clock,reset);
    assign seq_loop_intf_177.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state6;
    assign seq_loop_intf_177.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_177.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_177.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_177.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state3;
    assign seq_loop_intf_177.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_177.post_loop_state1 = 9'h0;
    assign seq_loop_intf_177.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_177.post_loop_state2 = 9'h0;
    assign seq_loop_intf_177.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_177.post_loop_state3 = 9'h0;
    assign seq_loop_intf_177.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_177.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state7;
    assign seq_loop_intf_177.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_177.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_177.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_177.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_CS_fsm;
    assign seq_loop_intf_177.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state7;
    assign seq_loop_intf_177.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state9;
    assign seq_loop_intf_177.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_177.iter_end_state1 = 9'h0;
    assign seq_loop_intf_177.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_177.one_state_loop = 1'b0;
    assign seq_loop_intf_177.one_state_block = 1'b0;
    assign seq_loop_intf_177.finish = finish;
    csv_file_dump seq_loop_csv_dumper_177;
    seq_loop_monitor #(9) seq_loop_monitor_177;
    seq_loop_intf#(9) seq_loop_intf_178(clock,reset);
    assign seq_loop_intf_178.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state2;
    assign seq_loop_intf_178.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_178.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_178.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_178.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state2;
    assign seq_loop_intf_178.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_178.post_loop_state1 = 9'h0;
    assign seq_loop_intf_178.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_178.post_loop_state2 = 9'h0;
    assign seq_loop_intf_178.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_178.post_loop_state3 = 9'h0;
    assign seq_loop_intf_178.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_178.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state3;
    assign seq_loop_intf_178.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_178.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_178.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_178.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_CS_fsm;
    assign seq_loop_intf_178.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state3;
    assign seq_loop_intf_178.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state7;
    assign seq_loop_intf_178.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_178.iter_end_state1 = 9'h0;
    assign seq_loop_intf_178.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_178.one_state_loop = 1'b0;
    assign seq_loop_intf_178.one_state_block = 1'b0;
    assign seq_loop_intf_178.finish = finish;
    csv_file_dump seq_loop_csv_dumper_178;
    seq_loop_monitor #(9) seq_loop_monitor_178;
    seq_loop_intf#(9) seq_loop_intf_179(clock,reset);
    assign seq_loop_intf_179.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state1;
    assign seq_loop_intf_179.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_179.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_179.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_179.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state1;
    assign seq_loop_intf_179.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_179.post_loop_state1 = 9'h0;
    assign seq_loop_intf_179.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_179.post_loop_state2 = 9'h0;
    assign seq_loop_intf_179.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_179.post_loop_state3 = 9'h0;
    assign seq_loop_intf_179.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_179.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state2;
    assign seq_loop_intf_179.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_179.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_179.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_179.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_CS_fsm;
    assign seq_loop_intf_179.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state2;
    assign seq_loop_intf_179.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_NTT2_ext_1_fu_3357.ap_ST_fsm_state3;
    assign seq_loop_intf_179.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_179.iter_end_state1 = 9'h0;
    assign seq_loop_intf_179.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_179.one_state_loop = 1'b0;
    assign seq_loop_intf_179.one_state_block = 1'b0;
    assign seq_loop_intf_179.finish = finish;
    csv_file_dump seq_loop_csv_dumper_179;
    seq_loop_monitor #(9) seq_loop_monitor_179;
    seq_loop_intf#(11) seq_loop_intf_180(clock,reset);
    assign seq_loop_intf_180.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state6;
    assign seq_loop_intf_180.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_180.pre_loop_state1 = 11'h0;
    assign seq_loop_intf_180.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_180.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state3;
    assign seq_loop_intf_180.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_180.post_loop_state1 = 11'h0;
    assign seq_loop_intf_180.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_180.post_loop_state2 = 11'h0;
    assign seq_loop_intf_180.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_180.post_loop_state3 = 11'h0;
    assign seq_loop_intf_180.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_180.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state7;
    assign seq_loop_intf_180.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_180.quit_loop_state1 = 11'h0;
    assign seq_loop_intf_180.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_180.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_CS_fsm;
    assign seq_loop_intf_180.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state7;
    assign seq_loop_intf_180.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state9;
    assign seq_loop_intf_180.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_180.iter_end_state1 = 11'h0;
    assign seq_loop_intf_180.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_180.one_state_loop = 1'b0;
    assign seq_loop_intf_180.one_state_block = 1'b0;
    assign seq_loop_intf_180.finish = finish;
    csv_file_dump seq_loop_csv_dumper_180;
    seq_loop_monitor #(11) seq_loop_monitor_180;
    seq_loop_intf#(11) seq_loop_intf_181(clock,reset);
    assign seq_loop_intf_181.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state2;
    assign seq_loop_intf_181.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_181.pre_loop_state1 = 11'h0;
    assign seq_loop_intf_181.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_181.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state2;
    assign seq_loop_intf_181.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_181.post_loop_state1 = 11'h0;
    assign seq_loop_intf_181.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_181.post_loop_state2 = 11'h0;
    assign seq_loop_intf_181.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_181.post_loop_state3 = 11'h0;
    assign seq_loop_intf_181.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_181.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state3;
    assign seq_loop_intf_181.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_181.quit_loop_state1 = 11'h0;
    assign seq_loop_intf_181.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_181.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_CS_fsm;
    assign seq_loop_intf_181.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state3;
    assign seq_loop_intf_181.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state7;
    assign seq_loop_intf_181.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_181.iter_end_state1 = 11'h0;
    assign seq_loop_intf_181.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_181.one_state_loop = 1'b0;
    assign seq_loop_intf_181.one_state_block = 1'b0;
    assign seq_loop_intf_181.finish = finish;
    csv_file_dump seq_loop_csv_dumper_181;
    seq_loop_monitor #(11) seq_loop_monitor_181;
    seq_loop_intf#(11) seq_loop_intf_182(clock,reset);
    assign seq_loop_intf_182.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state1;
    assign seq_loop_intf_182.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_182.pre_loop_state1 = 11'h0;
    assign seq_loop_intf_182.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_182.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state10;
    assign seq_loop_intf_182.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_182.post_loop_state1 = 11'h0;
    assign seq_loop_intf_182.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_182.post_loop_state2 = 11'h0;
    assign seq_loop_intf_182.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_182.post_loop_state3 = 11'h0;
    assign seq_loop_intf_182.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_182.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state2;
    assign seq_loop_intf_182.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_182.quit_loop_state1 = 11'h0;
    assign seq_loop_intf_182.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_182.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_CS_fsm;
    assign seq_loop_intf_182.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state2;
    assign seq_loop_intf_182.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state3;
    assign seq_loop_intf_182.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_182.iter_end_state1 = 11'h0;
    assign seq_loop_intf_182.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_182.one_state_loop = 1'b0;
    assign seq_loop_intf_182.one_state_block = 1'b0;
    assign seq_loop_intf_182.finish = finish;
    csv_file_dump seq_loop_csv_dumper_182;
    seq_loop_monitor #(11) seq_loop_monitor_182;
    seq_loop_intf#(11) seq_loop_intf_183(clock,reset);
    assign seq_loop_intf_183.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state1;
    assign seq_loop_intf_183.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_183.pre_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state2;
    assign seq_loop_intf_183.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_183.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state1;
    assign seq_loop_intf_183.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_183.post_loop_state1 = 11'h0;
    assign seq_loop_intf_183.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_183.post_loop_state2 = 11'h0;
    assign seq_loop_intf_183.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_183.post_loop_state3 = 11'h0;
    assign seq_loop_intf_183.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_183.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state10;
    assign seq_loop_intf_183.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_183.quit_loop_state1 = 11'h0;
    assign seq_loop_intf_183.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_183.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_CS_fsm;
    assign seq_loop_intf_183.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state10;
    assign seq_loop_intf_183.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_modp_iNTT2_ext_1_fu_3386.ap_ST_fsm_state11;
    assign seq_loop_intf_183.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_183.iter_end_state1 = 11'h0;
    assign seq_loop_intf_183.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_183.one_state_loop = 1'b0;
    assign seq_loop_intf_183.one_state_block = 1'b0;
    assign seq_loop_intf_183.finish = finish;
    csv_file_dump seq_loop_csv_dumper_183;
    seq_loop_monitor #(11) seq_loop_monitor_183;
    seq_loop_intf#(13) seq_loop_intf_184(clock,reset);
    assign seq_loop_intf_184.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state4;
    assign seq_loop_intf_184.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_184.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_184.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_184.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state3;
    assign seq_loop_intf_184.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_184.post_loop_state1 = 13'h0;
    assign seq_loop_intf_184.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_184.post_loop_state2 = 13'h0;
    assign seq_loop_intf_184.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_184.post_loop_state3 = 13'h0;
    assign seq_loop_intf_184.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_184.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state5;
    assign seq_loop_intf_184.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_184.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_184.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_184.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_CS_fsm;
    assign seq_loop_intf_184.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state5;
    assign seq_loop_intf_184.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state13;
    assign seq_loop_intf_184.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_184.iter_end_state1 = 13'h0;
    assign seq_loop_intf_184.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_184.one_state_loop = 1'b0;
    assign seq_loop_intf_184.one_state_block = 1'b0;
    assign seq_loop_intf_184.finish = finish;
    csv_file_dump seq_loop_csv_dumper_184;
    seq_loop_monitor #(13) seq_loop_monitor_184;
    seq_loop_intf#(13) seq_loop_intf_185(clock,reset);
    assign seq_loop_intf_185.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state2;
    assign seq_loop_intf_185.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_185.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_185.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_185.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state2;
    assign seq_loop_intf_185.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_185.post_loop_state1 = 13'h0;
    assign seq_loop_intf_185.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_185.post_loop_state2 = 13'h0;
    assign seq_loop_intf_185.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_185.post_loop_state3 = 13'h0;
    assign seq_loop_intf_185.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_185.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state3;
    assign seq_loop_intf_185.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_185.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_185.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_185.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_CS_fsm;
    assign seq_loop_intf_185.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state3;
    assign seq_loop_intf_185.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state5;
    assign seq_loop_intf_185.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_185.iter_end_state1 = 13'h0;
    assign seq_loop_intf_185.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_185.one_state_loop = 1'b0;
    assign seq_loop_intf_185.one_state_block = 1'b0;
    assign seq_loop_intf_185.finish = finish;
    csv_file_dump seq_loop_csv_dumper_185;
    seq_loop_monitor #(13) seq_loop_monitor_185;
    seq_loop_intf#(13) seq_loop_intf_186(clock,reset);
    assign seq_loop_intf_186.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state1;
    assign seq_loop_intf_186.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_186.pre_loop_state1 = 13'h0;
    assign seq_loop_intf_186.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_186.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state1;
    assign seq_loop_intf_186.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_186.post_loop_state1 = 13'h0;
    assign seq_loop_intf_186.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_186.post_loop_state2 = 13'h0;
    assign seq_loop_intf_186.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_186.post_loop_state3 = 13'h0;
    assign seq_loop_intf_186.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_186.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state2;
    assign seq_loop_intf_186.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_186.quit_loop_state1 = 13'h0;
    assign seq_loop_intf_186.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_186.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_CS_fsm;
    assign seq_loop_intf_186.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state2;
    assign seq_loop_intf_186.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_FFT_1_fu_3500.ap_ST_fsm_state3;
    assign seq_loop_intf_186.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_186.iter_end_state1 = 13'h0;
    assign seq_loop_intf_186.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_186.one_state_loop = 1'b0;
    assign seq_loop_intf_186.one_state_block = 1'b0;
    assign seq_loop_intf_186.finish = finish;
    csv_file_dump seq_loop_csv_dumper_186;
    seq_loop_monitor #(13) seq_loop_monitor_186;
    seq_loop_intf#(17) seq_loop_intf_187(clock,reset);
    assign seq_loop_intf_187.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state4;
    assign seq_loop_intf_187.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_187.pre_loop_state1 = 17'h0;
    assign seq_loop_intf_187.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_187.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state3;
    assign seq_loop_intf_187.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_187.post_loop_state1 = 17'h0;
    assign seq_loop_intf_187.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_187.post_loop_state2 = 17'h0;
    assign seq_loop_intf_187.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_187.post_loop_state3 = 17'h0;
    assign seq_loop_intf_187.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_187.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state5;
    assign seq_loop_intf_187.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_187.quit_loop_state1 = 17'h0;
    assign seq_loop_intf_187.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_187.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_CS_fsm;
    assign seq_loop_intf_187.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state5;
    assign seq_loop_intf_187.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state13;
    assign seq_loop_intf_187.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_187.iter_end_state1 = 17'h0;
    assign seq_loop_intf_187.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_187.one_state_loop = 1'b0;
    assign seq_loop_intf_187.one_state_block = 1'b0;
    assign seq_loop_intf_187.finish = finish;
    csv_file_dump seq_loop_csv_dumper_187;
    seq_loop_monitor #(17) seq_loop_monitor_187;
    seq_loop_intf#(17) seq_loop_intf_188(clock,reset);
    assign seq_loop_intf_188.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state2;
    assign seq_loop_intf_188.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_188.pre_loop_state1 = 17'h0;
    assign seq_loop_intf_188.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_188.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state2;
    assign seq_loop_intf_188.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_188.post_loop_state1 = 17'h0;
    assign seq_loop_intf_188.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_188.post_loop_state2 = 17'h0;
    assign seq_loop_intf_188.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_188.post_loop_state3 = 17'h0;
    assign seq_loop_intf_188.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_188.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state3;
    assign seq_loop_intf_188.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_188.quit_loop_state1 = 17'h0;
    assign seq_loop_intf_188.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_188.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_CS_fsm;
    assign seq_loop_intf_188.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state3;
    assign seq_loop_intf_188.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state5;
    assign seq_loop_intf_188.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_188.iter_end_state1 = 17'h0;
    assign seq_loop_intf_188.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_188.one_state_loop = 1'b0;
    assign seq_loop_intf_188.one_state_block = 1'b0;
    assign seq_loop_intf_188.finish = finish;
    csv_file_dump seq_loop_csv_dumper_188;
    seq_loop_monitor #(17) seq_loop_monitor_188;
    seq_loop_intf#(17) seq_loop_intf_189(clock,reset);
    assign seq_loop_intf_189.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state1;
    assign seq_loop_intf_189.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_189.pre_loop_state1 = 17'h0;
    assign seq_loop_intf_189.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_189.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state14;
    assign seq_loop_intf_189.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_189.post_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state15;
    assign seq_loop_intf_189.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_189.post_loop_state2 = 17'h0;
    assign seq_loop_intf_189.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_189.post_loop_state3 = 17'h0;
    assign seq_loop_intf_189.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_189.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state2;
    assign seq_loop_intf_189.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_189.quit_loop_state1 = 17'h0;
    assign seq_loop_intf_189.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_189.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_CS_fsm;
    assign seq_loop_intf_189.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state2;
    assign seq_loop_intf_189.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state3;
    assign seq_loop_intf_189.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_189.iter_end_state1 = 17'h0;
    assign seq_loop_intf_189.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_189.one_state_loop = 1'b0;
    assign seq_loop_intf_189.one_state_block = 1'b0;
    assign seq_loop_intf_189.finish = finish;
    csv_file_dump seq_loop_csv_dumper_189;
    seq_loop_monitor #(17) seq_loop_monitor_189;
    seq_loop_intf#(17) seq_loop_intf_190(clock,reset);
    assign seq_loop_intf_190.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state2;
    assign seq_loop_intf_190.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_190.pre_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state14;
    assign seq_loop_intf_190.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_190.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state1;
    assign seq_loop_intf_190.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_190.post_loop_state1 = 17'h0;
    assign seq_loop_intf_190.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_190.post_loop_state2 = 17'h0;
    assign seq_loop_intf_190.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_190.post_loop_state3 = 17'h0;
    assign seq_loop_intf_190.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_190.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state15;
    assign seq_loop_intf_190.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_190.quit_loop_state1 = 17'h0;
    assign seq_loop_intf_190.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_190.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_CS_fsm;
    assign seq_loop_intf_190.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state15;
    assign seq_loop_intf_190.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_iFFT_1_fu_3522.ap_ST_fsm_state17;
    assign seq_loop_intf_190.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_190.iter_end_state1 = 17'h0;
    assign seq_loop_intf_190.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_190.one_state_loop = 1'b0;
    assign seq_loop_intf_190.one_state_block = 1'b0;
    assign seq_loop_intf_190.finish = finish;
    csv_file_dump seq_loop_csv_dumper_190;
    seq_loop_monitor #(17) seq_loop_monitor_190;
    seq_loop_intf#(4) seq_loop_intf_191(clock,reset);
    assign seq_loop_intf_191.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_mod_small_signed_1_fu_3545.ap_ST_fsm_state1;
    assign seq_loop_intf_191.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_191.pre_loop_state1 = 4'h0;
    assign seq_loop_intf_191.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_191.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_mod_small_signed_1_fu_3545.ap_ST_fsm_state4;
    assign seq_loop_intf_191.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_191.post_loop_state1 = 4'h0;
    assign seq_loop_intf_191.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_191.post_loop_state2 = 4'h0;
    assign seq_loop_intf_191.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_191.post_loop_state3 = 4'h0;
    assign seq_loop_intf_191.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_191.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_mod_small_signed_1_fu_3545.ap_ST_fsm_state3;
    assign seq_loop_intf_191.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_191.quit_loop_state1 = 4'h0;
    assign seq_loop_intf_191.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_191.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_mod_small_signed_1_fu_3545.ap_CS_fsm;
    assign seq_loop_intf_191.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_mod_small_signed_1_fu_3545.ap_ST_fsm_state2;
    assign seq_loop_intf_191.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_mod_small_signed_1_fu_3545.ap_ST_fsm_state3;
    assign seq_loop_intf_191.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_191.iter_end_state1 = 4'h0;
    assign seq_loop_intf_191.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_191.one_state_loop = 1'b0;
    assign seq_loop_intf_191.one_state_block = 1'b0;
    assign seq_loop_intf_191.finish = finish;
    csv_file_dump seq_loop_csv_dumper_191;
    seq_loop_monitor #(4) seq_loop_monitor_191;
    seq_loop_intf#(19) seq_loop_intf_192(clock,reset);
    assign seq_loop_intf_192.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state8;
    assign seq_loop_intf_192.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_192.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_192.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_192.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state11;
    assign seq_loop_intf_192.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_192.post_loop_state1 = 19'h0;
    assign seq_loop_intf_192.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_192.post_loop_state2 = 19'h0;
    assign seq_loop_intf_192.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_192.post_loop_state3 = 19'h0;
    assign seq_loop_intf_192.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_192.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state10;
    assign seq_loop_intf_192.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_192.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_192.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_192.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_CS_fsm;
    assign seq_loop_intf_192.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state9;
    assign seq_loop_intf_192.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state10;
    assign seq_loop_intf_192.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_192.iter_end_state1 = 19'h0;
    assign seq_loop_intf_192.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_192.one_state_loop = 1'b0;
    assign seq_loop_intf_192.one_state_block = 1'b0;
    assign seq_loop_intf_192.finish = finish;
    csv_file_dump seq_loop_csv_dumper_192;
    seq_loop_monitor #(19) seq_loop_monitor_192;
    seq_loop_intf#(19) seq_loop_intf_193(clock,reset);
    assign seq_loop_intf_193.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state10;
    assign seq_loop_intf_193.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_193.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_193.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_193.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state7;
    assign seq_loop_intf_193.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_193.post_loop_state1 = 19'h0;
    assign seq_loop_intf_193.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_193.post_loop_state2 = 19'h0;
    assign seq_loop_intf_193.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_193.post_loop_state3 = 19'h0;
    assign seq_loop_intf_193.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_193.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state11;
    assign seq_loop_intf_193.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_193.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_193.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_193.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_CS_fsm;
    assign seq_loop_intf_193.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state11;
    assign seq_loop_intf_193.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state12;
    assign seq_loop_intf_193.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_193.iter_end_state1 = 19'h0;
    assign seq_loop_intf_193.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_193.one_state_loop = 1'b0;
    assign seq_loop_intf_193.one_state_block = 1'b0;
    assign seq_loop_intf_193.finish = finish;
    csv_file_dump seq_loop_csv_dumper_193;
    seq_loop_monitor #(19) seq_loop_monitor_193;
    seq_loop_intf#(19) seq_loop_intf_194(clock,reset);
    assign seq_loop_intf_194.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state6;
    assign seq_loop_intf_194.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_194.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_194.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_194.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state13;
    assign seq_loop_intf_194.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_194.post_loop_state1 = 19'h0;
    assign seq_loop_intf_194.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_194.post_loop_state2 = 19'h0;
    assign seq_loop_intf_194.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_194.post_loop_state3 = 19'h0;
    assign seq_loop_intf_194.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_194.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state7;
    assign seq_loop_intf_194.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_194.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_194.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_194.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_CS_fsm;
    assign seq_loop_intf_194.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state7;
    assign seq_loop_intf_194.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state11;
    assign seq_loop_intf_194.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_194.iter_end_state1 = 19'h0;
    assign seq_loop_intf_194.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_194.one_state_loop = 1'b0;
    assign seq_loop_intf_194.one_state_block = 1'b0;
    assign seq_loop_intf_194.finish = finish;
    csv_file_dump seq_loop_csv_dumper_194;
    seq_loop_monitor #(19) seq_loop_monitor_194;
    seq_loop_intf#(19) seq_loop_intf_195(clock,reset);
    assign seq_loop_intf_195.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state7;
    assign seq_loop_intf_195.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_195.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_195.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_195.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state2;
    assign seq_loop_intf_195.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_195.post_loop_state1 = 19'h0;
    assign seq_loop_intf_195.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_195.post_loop_state2 = 19'h0;
    assign seq_loop_intf_195.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_195.post_loop_state3 = 19'h0;
    assign seq_loop_intf_195.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_195.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state13;
    assign seq_loop_intf_195.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_195.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_195.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_195.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_CS_fsm;
    assign seq_loop_intf_195.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state13;
    assign seq_loop_intf_195.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state14;
    assign seq_loop_intf_195.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_195.iter_end_state1 = 19'h0;
    assign seq_loop_intf_195.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_195.one_state_loop = 1'b0;
    assign seq_loop_intf_195.one_state_block = 1'b0;
    assign seq_loop_intf_195.finish = finish;
    csv_file_dump seq_loop_csv_dumper_195;
    seq_loop_monitor #(19) seq_loop_monitor_195;
    seq_loop_intf#(19) seq_loop_intf_196(clock,reset);
    assign seq_loop_intf_196.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state1;
    assign seq_loop_intf_196.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_196.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_196.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_196.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state15;
    assign seq_loop_intf_196.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_196.post_loop_state1 = 19'h0;
    assign seq_loop_intf_196.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_196.post_loop_state2 = 19'h0;
    assign seq_loop_intf_196.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_196.post_loop_state3 = 19'h0;
    assign seq_loop_intf_196.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_196.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state2;
    assign seq_loop_intf_196.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_196.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_196.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_196.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_CS_fsm;
    assign seq_loop_intf_196.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state2;
    assign seq_loop_intf_196.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state13;
    assign seq_loop_intf_196.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_196.iter_end_state1 = 19'h0;
    assign seq_loop_intf_196.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_196.one_state_loop = 1'b0;
    assign seq_loop_intf_196.one_state_block = 1'b0;
    assign seq_loop_intf_196.finish = finish;
    csv_file_dump seq_loop_csv_dumper_196;
    seq_loop_monitor #(19) seq_loop_monitor_196;
    seq_loop_intf#(19) seq_loop_intf_197(clock,reset);
    assign seq_loop_intf_197.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state15;
    assign seq_loop_intf_197.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_197.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_197.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_197.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state18;
    assign seq_loop_intf_197.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_197.post_loop_state1 = 19'h0;
    assign seq_loop_intf_197.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_197.post_loop_state2 = 19'h0;
    assign seq_loop_intf_197.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_197.post_loop_state3 = 19'h0;
    assign seq_loop_intf_197.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_197.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state17;
    assign seq_loop_intf_197.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_197.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_197.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_197.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_CS_fsm;
    assign seq_loop_intf_197.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state16;
    assign seq_loop_intf_197.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state17;
    assign seq_loop_intf_197.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_197.iter_end_state1 = 19'h0;
    assign seq_loop_intf_197.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_197.one_state_loop = 1'b0;
    assign seq_loop_intf_197.one_state_block = 1'b0;
    assign seq_loop_intf_197.finish = finish;
    csv_file_dump seq_loop_csv_dumper_197;
    seq_loop_monitor #(19) seq_loop_monitor_197;
    seq_loop_intf#(19) seq_loop_intf_198(clock,reset);
    assign seq_loop_intf_198.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state17;
    assign seq_loop_intf_198.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_198.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_198.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_198.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state15;
    assign seq_loop_intf_198.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_198.post_loop_state1 = 19'h0;
    assign seq_loop_intf_198.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_198.post_loop_state2 = 19'h0;
    assign seq_loop_intf_198.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_198.post_loop_state3 = 19'h0;
    assign seq_loop_intf_198.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_198.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state18;
    assign seq_loop_intf_198.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_198.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_198.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_198.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_CS_fsm;
    assign seq_loop_intf_198.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state18;
    assign seq_loop_intf_198.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state19;
    assign seq_loop_intf_198.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_198.iter_end_state1 = 19'h0;
    assign seq_loop_intf_198.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_198.one_state_loop = 1'b0;
    assign seq_loop_intf_198.one_state_block = 1'b0;
    assign seq_loop_intf_198.finish = finish;
    csv_file_dump seq_loop_csv_dumper_198;
    seq_loop_monitor #(19) seq_loop_monitor_198;
    seq_loop_intf#(19) seq_loop_intf_199(clock,reset);
    assign seq_loop_intf_199.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state2;
    assign seq_loop_intf_199.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_199.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_199.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_199.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state1;
    assign seq_loop_intf_199.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_199.post_loop_state1 = 19'h0;
    assign seq_loop_intf_199.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_199.post_loop_state2 = 19'h0;
    assign seq_loop_intf_199.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_199.post_loop_state3 = 19'h0;
    assign seq_loop_intf_199.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_199.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state15;
    assign seq_loop_intf_199.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_199.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_199.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_199.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_CS_fsm;
    assign seq_loop_intf_199.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state15;
    assign seq_loop_intf_199.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_rebuild_CRT_1_fu_3561.ap_ST_fsm_state18;
    assign seq_loop_intf_199.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_199.iter_end_state1 = 19'h0;
    assign seq_loop_intf_199.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_199.one_state_loop = 1'b0;
    assign seq_loop_intf_199.one_state_block = 1'b0;
    assign seq_loop_intf_199.finish = finish;
    csv_file_dump seq_loop_csv_dumper_199;
    seq_loop_monitor #(19) seq_loop_monitor_199;
    seq_loop_intf#(8) seq_loop_intf_200(clock,reset);
    assign seq_loop_intf_200.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state1;
    assign seq_loop_intf_200.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_200.pre_loop_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state4;
    assign seq_loop_intf_200.pre_states_valid[1] = 1'b1;
    assign seq_loop_intf_200.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state3;
    assign seq_loop_intf_200.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_200.post_loop_state1 = 8'h0;
    assign seq_loop_intf_200.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_200.post_loop_state2 = 8'h0;
    assign seq_loop_intf_200.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_200.post_loop_state3 = 8'h0;
    assign seq_loop_intf_200.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_200.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state2;
    assign seq_loop_intf_200.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_200.quit_loop_state1 = 8'h0;
    assign seq_loop_intf_200.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_200.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_CS_fsm;
    assign seq_loop_intf_200.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state2;
    assign seq_loop_intf_200.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state2;
    assign seq_loop_intf_200.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_200.iter_end_state1 = 8'h0;
    assign seq_loop_intf_200.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_200.one_state_loop = 1'b1;
    assign seq_loop_intf_200.one_state_block = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state2_blk;
    assign seq_loop_intf_200.finish = finish;
    csv_file_dump seq_loop_csv_dumper_200;
    seq_loop_monitor #(8) seq_loop_monitor_200;
    seq_loop_intf#(8) seq_loop_intf_201(clock,reset);
    assign seq_loop_intf_201.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state3;
    assign seq_loop_intf_201.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_201.pre_loop_state1 = 8'h0;
    assign seq_loop_intf_201.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_201.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state2;
    assign seq_loop_intf_201.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_201.post_loop_state1 = 8'h0;
    assign seq_loop_intf_201.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_201.post_loop_state2 = 8'h0;
    assign seq_loop_intf_201.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_201.post_loop_state3 = 8'h0;
    assign seq_loop_intf_201.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_201.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state4;
    assign seq_loop_intf_201.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_201.quit_loop_state1 = 8'h0;
    assign seq_loop_intf_201.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_201.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_CS_fsm;
    assign seq_loop_intf_201.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state4;
    assign seq_loop_intf_201.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state8;
    assign seq_loop_intf_201.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_201.iter_end_state1 = 8'h0;
    assign seq_loop_intf_201.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_201.one_state_loop = 1'b0;
    assign seq_loop_intf_201.one_state_block = 1'b0;
    assign seq_loop_intf_201.finish = finish;
    csv_file_dump seq_loop_csv_dumper_201;
    seq_loop_monitor #(8) seq_loop_monitor_201;
    seq_loop_intf#(8) seq_loop_intf_202(clock,reset);
    assign seq_loop_intf_202.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state1;
    assign seq_loop_intf_202.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_202.pre_loop_state1 = 8'h0;
    assign seq_loop_intf_202.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_202.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state1;
    assign seq_loop_intf_202.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_202.post_loop_state1 = 8'h0;
    assign seq_loop_intf_202.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_202.post_loop_state2 = 8'h0;
    assign seq_loop_intf_202.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_202.post_loop_state3 = 8'h0;
    assign seq_loop_intf_202.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_202.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state2;
    assign seq_loop_intf_202.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_202.quit_loop_state1 = 8'h0;
    assign seq_loop_intf_202.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_202.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_CS_fsm;
    assign seq_loop_intf_202.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state2;
    assign seq_loop_intf_202.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state4;
    assign seq_loop_intf_202.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_202.iter_end_state1 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_big_to_fp_1_fu_3592.ap_ST_fsm_state2;
    assign seq_loop_intf_202.iter_end_states_valid[1] = 1'b1;
    assign seq_loop_intf_202.one_state_loop = 1'b0;
    assign seq_loop_intf_202.one_state_block = 1'b0;
    assign seq_loop_intf_202.finish = finish;
    csv_file_dump seq_loop_csv_dumper_202;
    seq_loop_monitor #(8) seq_loop_monitor_202;
    seq_loop_intf#(9) seq_loop_intf_203(clock,reset);
    assign seq_loop_intf_203.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_mul_fft_1_fu_3613.ap_ST_fsm_state1;
    assign seq_loop_intf_203.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_203.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_203.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_203.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_mul_fft_1_fu_3613.ap_ST_fsm_state1;
    assign seq_loop_intf_203.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_203.post_loop_state1 = 9'h0;
    assign seq_loop_intf_203.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_203.post_loop_state2 = 9'h0;
    assign seq_loop_intf_203.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_203.post_loop_state3 = 9'h0;
    assign seq_loop_intf_203.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_203.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_mul_fft_1_fu_3613.ap_ST_fsm_state2;
    assign seq_loop_intf_203.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_203.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_203.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_203.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_mul_fft_1_fu_3613.ap_CS_fsm;
    assign seq_loop_intf_203.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_mul_fft_1_fu_3613.ap_ST_fsm_state2;
    assign seq_loop_intf_203.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_mul_fft_1_fu_3613.ap_ST_fsm_state9;
    assign seq_loop_intf_203.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_203.iter_end_state1 = 9'h0;
    assign seq_loop_intf_203.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_203.one_state_loop = 1'b0;
    assign seq_loop_intf_203.one_state_block = 1'b0;
    assign seq_loop_intf_203.finish = finish;
    csv_file_dump seq_loop_csv_dumper_203;
    seq_loop_monitor #(9) seq_loop_monitor_203;
    seq_loop_intf#(33) seq_loop_intf_204(clock,reset);
    assign seq_loop_intf_204.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state2;
    assign seq_loop_intf_204.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_204.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_204.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_204.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state5;
    assign seq_loop_intf_204.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_204.post_loop_state1 = 33'h0;
    assign seq_loop_intf_204.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_204.post_loop_state2 = 33'h0;
    assign seq_loop_intf_204.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_204.post_loop_state3 = 33'h0;
    assign seq_loop_intf_204.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_204.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state4;
    assign seq_loop_intf_204.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_204.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_204.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_204.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_204.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state3;
    assign seq_loop_intf_204.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state4;
    assign seq_loop_intf_204.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_204.iter_end_state1 = 33'h0;
    assign seq_loop_intf_204.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_204.one_state_loop = 1'b0;
    assign seq_loop_intf_204.one_state_block = 1'b0;
    assign seq_loop_intf_204.finish = finish;
    csv_file_dump seq_loop_csv_dumper_204;
    seq_loop_monitor #(33) seq_loop_monitor_204;
    seq_loop_intf#(33) seq_loop_intf_205(clock,reset);
    assign seq_loop_intf_205.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state4;
    assign seq_loop_intf_205.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_205.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_205.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_205.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state7;
    assign seq_loop_intf_205.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_205.post_loop_state1 = 33'h0;
    assign seq_loop_intf_205.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_205.post_loop_state2 = 33'h0;
    assign seq_loop_intf_205.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_205.post_loop_state3 = 33'h0;
    assign seq_loop_intf_205.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_205.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state6;
    assign seq_loop_intf_205.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_205.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_205.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_205.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_205.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state5;
    assign seq_loop_intf_205.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state6;
    assign seq_loop_intf_205.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_205.iter_end_state1 = 33'h0;
    assign seq_loop_intf_205.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_205.one_state_loop = 1'b0;
    assign seq_loop_intf_205.one_state_block = 1'b0;
    assign seq_loop_intf_205.finish = finish;
    csv_file_dump seq_loop_csv_dumper_205;
    seq_loop_monitor #(33) seq_loop_monitor_205;
    seq_loop_intf#(33) seq_loop_intf_206(clock,reset);
    assign seq_loop_intf_206.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state7;
    assign seq_loop_intf_206.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_206.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_206.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_206.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state9;
    assign seq_loop_intf_206.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_206.post_loop_state1 = 33'h0;
    assign seq_loop_intf_206.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_206.post_loop_state2 = 33'h0;
    assign seq_loop_intf_206.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_206.post_loop_state3 = 33'h0;
    assign seq_loop_intf_206.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_206.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state8;
    assign seq_loop_intf_206.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_206.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_206.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_206.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_206.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state8;
    assign seq_loop_intf_206.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state8;
    assign seq_loop_intf_206.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_206.iter_end_state1 = 33'h0;
    assign seq_loop_intf_206.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_206.one_state_loop = 1'b1;
    assign seq_loop_intf_206.one_state_block = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state8_blk;
    assign seq_loop_intf_206.finish = finish;
    csv_file_dump seq_loop_csv_dumper_206;
    seq_loop_monitor #(33) seq_loop_monitor_206;
    seq_loop_intf#(33) seq_loop_intf_207(clock,reset);
    assign seq_loop_intf_207.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state8;
    assign seq_loop_intf_207.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_207.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_207.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_207.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state10;
    assign seq_loop_intf_207.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_207.post_loop_state1 = 33'h0;
    assign seq_loop_intf_207.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_207.post_loop_state2 = 33'h0;
    assign seq_loop_intf_207.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_207.post_loop_state3 = 33'h0;
    assign seq_loop_intf_207.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_207.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state9;
    assign seq_loop_intf_207.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_207.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_207.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_207.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_207.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state9;
    assign seq_loop_intf_207.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state9;
    assign seq_loop_intf_207.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_207.iter_end_state1 = 33'h0;
    assign seq_loop_intf_207.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_207.one_state_loop = 1'b1;
    assign seq_loop_intf_207.one_state_block = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state9_blk;
    assign seq_loop_intf_207.finish = finish;
    csv_file_dump seq_loop_csv_dumper_207;
    seq_loop_monitor #(33) seq_loop_monitor_207;
    seq_loop_intf#(33) seq_loop_intf_208(clock,reset);
    assign seq_loop_intf_208.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state9;
    assign seq_loop_intf_208.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_208.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_208.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_208.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state12;
    assign seq_loop_intf_208.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_208.post_loop_state1 = 33'h0;
    assign seq_loop_intf_208.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_208.post_loop_state2 = 33'h0;
    assign seq_loop_intf_208.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_208.post_loop_state3 = 33'h0;
    assign seq_loop_intf_208.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_208.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state11;
    assign seq_loop_intf_208.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_208.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_208.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_208.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_208.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state10;
    assign seq_loop_intf_208.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state11;
    assign seq_loop_intf_208.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_208.iter_end_state1 = 33'h0;
    assign seq_loop_intf_208.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_208.one_state_loop = 1'b0;
    assign seq_loop_intf_208.one_state_block = 1'b0;
    assign seq_loop_intf_208.finish = finish;
    csv_file_dump seq_loop_csv_dumper_208;
    seq_loop_monitor #(33) seq_loop_monitor_208;
    seq_loop_intf#(33) seq_loop_intf_209(clock,reset);
    assign seq_loop_intf_209.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state11;
    assign seq_loop_intf_209.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_209.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_209.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_209.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state14;
    assign seq_loop_intf_209.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_209.post_loop_state1 = 33'h0;
    assign seq_loop_intf_209.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_209.post_loop_state2 = 33'h0;
    assign seq_loop_intf_209.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_209.post_loop_state3 = 33'h0;
    assign seq_loop_intf_209.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_209.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state13;
    assign seq_loop_intf_209.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_209.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_209.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_209.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_209.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state12;
    assign seq_loop_intf_209.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state13;
    assign seq_loop_intf_209.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_209.iter_end_state1 = 33'h0;
    assign seq_loop_intf_209.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_209.one_state_loop = 1'b0;
    assign seq_loop_intf_209.one_state_block = 1'b0;
    assign seq_loop_intf_209.finish = finish;
    csv_file_dump seq_loop_csv_dumper_209;
    seq_loop_monitor #(33) seq_loop_monitor_209;
    seq_loop_intf#(33) seq_loop_intf_210(clock,reset);
    assign seq_loop_intf_210.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state16;
    assign seq_loop_intf_210.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_210.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_210.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_210.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state19;
    assign seq_loop_intf_210.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_210.post_loop_state1 = 33'h0;
    assign seq_loop_intf_210.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_210.post_loop_state2 = 33'h0;
    assign seq_loop_intf_210.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_210.post_loop_state3 = 33'h0;
    assign seq_loop_intf_210.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_210.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state18;
    assign seq_loop_intf_210.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_210.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_210.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_210.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_210.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state17;
    assign seq_loop_intf_210.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state18;
    assign seq_loop_intf_210.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_210.iter_end_state1 = 33'h0;
    assign seq_loop_intf_210.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_210.one_state_loop = 1'b0;
    assign seq_loop_intf_210.one_state_block = 1'b0;
    assign seq_loop_intf_210.finish = finish;
    csv_file_dump seq_loop_csv_dumper_210;
    seq_loop_monitor #(33) seq_loop_monitor_210;
    seq_loop_intf#(33) seq_loop_intf_211(clock,reset);
    assign seq_loop_intf_211.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state19;
    assign seq_loop_intf_211.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_211.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_211.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_211.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state21;
    assign seq_loop_intf_211.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_211.post_loop_state1 = 33'h0;
    assign seq_loop_intf_211.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_211.post_loop_state2 = 33'h0;
    assign seq_loop_intf_211.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_211.post_loop_state3 = 33'h0;
    assign seq_loop_intf_211.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_211.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state20;
    assign seq_loop_intf_211.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_211.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_211.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_211.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_211.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state20;
    assign seq_loop_intf_211.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state20;
    assign seq_loop_intf_211.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_211.iter_end_state1 = 33'h0;
    assign seq_loop_intf_211.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_211.one_state_loop = 1'b1;
    assign seq_loop_intf_211.one_state_block = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state20_blk;
    assign seq_loop_intf_211.finish = finish;
    csv_file_dump seq_loop_csv_dumper_211;
    seq_loop_monitor #(33) seq_loop_monitor_211;
    seq_loop_intf#(33) seq_loop_intf_212(clock,reset);
    assign seq_loop_intf_212.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state20;
    assign seq_loop_intf_212.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_212.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_212.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_212.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state23;
    assign seq_loop_intf_212.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_212.post_loop_state1 = 33'h0;
    assign seq_loop_intf_212.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_212.post_loop_state2 = 33'h0;
    assign seq_loop_intf_212.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_212.post_loop_state3 = 33'h0;
    assign seq_loop_intf_212.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_212.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state21;
    assign seq_loop_intf_212.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_212.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_212.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_212.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_212.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state21;
    assign seq_loop_intf_212.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state22;
    assign seq_loop_intf_212.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_212.iter_end_state1 = 33'h0;
    assign seq_loop_intf_212.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_212.one_state_loop = 1'b0;
    assign seq_loop_intf_212.one_state_block = 1'b0;
    assign seq_loop_intf_212.finish = finish;
    csv_file_dump seq_loop_csv_dumper_212;
    seq_loop_monitor #(33) seq_loop_monitor_212;
    seq_loop_intf#(33) seq_loop_intf_213(clock,reset);
    assign seq_loop_intf_213.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state21;
    assign seq_loop_intf_213.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_213.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_213.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_213.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state25;
    assign seq_loop_intf_213.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_213.post_loop_state1 = 33'h0;
    assign seq_loop_intf_213.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_213.post_loop_state2 = 33'h0;
    assign seq_loop_intf_213.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_213.post_loop_state3 = 33'h0;
    assign seq_loop_intf_213.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_213.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state23;
    assign seq_loop_intf_213.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_213.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_213.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_213.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_213.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state23;
    assign seq_loop_intf_213.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state24;
    assign seq_loop_intf_213.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_213.iter_end_state1 = 33'h0;
    assign seq_loop_intf_213.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_213.one_state_loop = 1'b0;
    assign seq_loop_intf_213.one_state_block = 1'b0;
    assign seq_loop_intf_213.finish = finish;
    csv_file_dump seq_loop_csv_dumper_213;
    seq_loop_monitor #(33) seq_loop_monitor_213;
    seq_loop_intf#(33) seq_loop_intf_214(clock,reset);
    assign seq_loop_intf_214.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state23;
    assign seq_loop_intf_214.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_214.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_214.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_214.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state27;
    assign seq_loop_intf_214.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_214.post_loop_state1 = 33'h0;
    assign seq_loop_intf_214.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_214.post_loop_state2 = 33'h0;
    assign seq_loop_intf_214.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_214.post_loop_state3 = 33'h0;
    assign seq_loop_intf_214.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_214.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state25;
    assign seq_loop_intf_214.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_214.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_214.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_214.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_214.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state25;
    assign seq_loop_intf_214.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state26;
    assign seq_loop_intf_214.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_214.iter_end_state1 = 33'h0;
    assign seq_loop_intf_214.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_214.one_state_loop = 1'b0;
    assign seq_loop_intf_214.one_state_block = 1'b0;
    assign seq_loop_intf_214.finish = finish;
    csv_file_dump seq_loop_csv_dumper_214;
    seq_loop_monitor #(33) seq_loop_monitor_214;
    seq_loop_intf#(33) seq_loop_intf_215(clock,reset);
    assign seq_loop_intf_215.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state15;
    assign seq_loop_intf_215.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_215.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_215.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_215.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state30;
    assign seq_loop_intf_215.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_215.post_loop_state1 = 33'h0;
    assign seq_loop_intf_215.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_215.post_loop_state2 = 33'h0;
    assign seq_loop_intf_215.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_215.post_loop_state3 = 33'h0;
    assign seq_loop_intf_215.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_215.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state16;
    assign seq_loop_intf_215.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_215.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_215.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_215.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_215.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state16;
    assign seq_loop_intf_215.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state29;
    assign seq_loop_intf_215.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_215.iter_end_state1 = 33'h0;
    assign seq_loop_intf_215.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_215.one_state_loop = 1'b0;
    assign seq_loop_intf_215.one_state_block = 1'b0;
    assign seq_loop_intf_215.finish = finish;
    csv_file_dump seq_loop_csv_dumper_215;
    seq_loop_monitor #(33) seq_loop_monitor_215;
    seq_loop_intf#(33) seq_loop_intf_216(clock,reset);
    assign seq_loop_intf_216.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state30;
    assign seq_loop_intf_216.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_216.pre_loop_state1 = 33'h0;
    assign seq_loop_intf_216.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_216.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state33;
    assign seq_loop_intf_216.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_216.post_loop_state1 = 33'h0;
    assign seq_loop_intf_216.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_216.post_loop_state2 = 33'h0;
    assign seq_loop_intf_216.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_216.post_loop_state3 = 33'h0;
    assign seq_loop_intf_216.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_216.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state31;
    assign seq_loop_intf_216.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_216.quit_loop_state1 = 33'h0;
    assign seq_loop_intf_216.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_216.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_CS_fsm;
    assign seq_loop_intf_216.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state31;
    assign seq_loop_intf_216.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.ap_ST_fsm_state32;
    assign seq_loop_intf_216.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_216.iter_end_state1 = 33'h0;
    assign seq_loop_intf_216.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_216.one_state_loop = 1'b0;
    assign seq_loop_intf_216.one_state_block = 1'b0;
    assign seq_loop_intf_216.finish = finish;
    csv_file_dump seq_loop_csv_dumper_216;
    seq_loop_monitor #(33) seq_loop_monitor_216;
    seq_loop_intf#(15) seq_loop_intf_217(clock,reset);
    assign seq_loop_intf_217.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state2;
    assign seq_loop_intf_217.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_217.pre_loop_state1 = 15'h0;
    assign seq_loop_intf_217.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_217.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state7;
    assign seq_loop_intf_217.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_217.post_loop_state1 = 15'h0;
    assign seq_loop_intf_217.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_217.post_loop_state2 = 15'h0;
    assign seq_loop_intf_217.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_217.post_loop_state3 = 15'h0;
    assign seq_loop_intf_217.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_217.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state3;
    assign seq_loop_intf_217.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_217.quit_loop_state1 = 15'h0;
    assign seq_loop_intf_217.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_217.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_CS_fsm;
    assign seq_loop_intf_217.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state3;
    assign seq_loop_intf_217.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state6;
    assign seq_loop_intf_217.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_217.iter_end_state1 = 15'h0;
    assign seq_loop_intf_217.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_217.one_state_loop = 1'b0;
    assign seq_loop_intf_217.one_state_block = 1'b0;
    assign seq_loop_intf_217.finish = finish;
    csv_file_dump seq_loop_csv_dumper_217;
    seq_loop_monitor #(15) seq_loop_monitor_217;
    seq_loop_intf#(15) seq_loop_intf_218(clock,reset);
    assign seq_loop_intf_218.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state7;
    assign seq_loop_intf_218.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_218.pre_loop_state1 = 15'h0;
    assign seq_loop_intf_218.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_218.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state10;
    assign seq_loop_intf_218.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_218.post_loop_state1 = 15'h0;
    assign seq_loop_intf_218.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_218.post_loop_state2 = 15'h0;
    assign seq_loop_intf_218.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_218.post_loop_state3 = 15'h0;
    assign seq_loop_intf_218.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_218.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state8;
    assign seq_loop_intf_218.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_218.quit_loop_state1 = 15'h0;
    assign seq_loop_intf_218.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_218.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_CS_fsm;
    assign seq_loop_intf_218.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state8;
    assign seq_loop_intf_218.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state9;
    assign seq_loop_intf_218.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_218.iter_end_state1 = 15'h0;
    assign seq_loop_intf_218.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_218.one_state_loop = 1'b0;
    assign seq_loop_intf_218.one_state_block = 1'b0;
    assign seq_loop_intf_218.finish = finish;
    csv_file_dump seq_loop_csv_dumper_218;
    seq_loop_monitor #(15) seq_loop_monitor_218;
    seq_loop_intf#(15) seq_loop_intf_219(clock,reset);
    assign seq_loop_intf_219.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state8;
    assign seq_loop_intf_219.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_219.pre_loop_state1 = 15'h0;
    assign seq_loop_intf_219.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_219.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state12;
    assign seq_loop_intf_219.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_219.post_loop_state1 = 15'h0;
    assign seq_loop_intf_219.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_219.post_loop_state2 = 15'h0;
    assign seq_loop_intf_219.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_219.post_loop_state3 = 15'h0;
    assign seq_loop_intf_219.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_219.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state10;
    assign seq_loop_intf_219.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_219.quit_loop_state1 = 15'h0;
    assign seq_loop_intf_219.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_219.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_CS_fsm;
    assign seq_loop_intf_219.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state10;
    assign seq_loop_intf_219.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state11;
    assign seq_loop_intf_219.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_219.iter_end_state1 = 15'h0;
    assign seq_loop_intf_219.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_219.one_state_loop = 1'b0;
    assign seq_loop_intf_219.one_state_block = 1'b0;
    assign seq_loop_intf_219.finish = finish;
    csv_file_dump seq_loop_csv_dumper_219;
    seq_loop_monitor #(15) seq_loop_monitor_219;
    seq_loop_intf#(15) seq_loop_intf_220(clock,reset);
    assign seq_loop_intf_220.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state10;
    assign seq_loop_intf_220.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_220.pre_loop_state1 = 15'h0;
    assign seq_loop_intf_220.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_220.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state14;
    assign seq_loop_intf_220.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_220.post_loop_state1 = 15'h0;
    assign seq_loop_intf_220.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_220.post_loop_state2 = 15'h0;
    assign seq_loop_intf_220.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_220.post_loop_state3 = 15'h0;
    assign seq_loop_intf_220.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_220.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state12;
    assign seq_loop_intf_220.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_220.quit_loop_state1 = 15'h0;
    assign seq_loop_intf_220.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_220.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_CS_fsm;
    assign seq_loop_intf_220.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state12;
    assign seq_loop_intf_220.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state13;
    assign seq_loop_intf_220.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_220.iter_end_state1 = 15'h0;
    assign seq_loop_intf_220.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_220.one_state_loop = 1'b0;
    assign seq_loop_intf_220.one_state_block = 1'b0;
    assign seq_loop_intf_220.finish = finish;
    csv_file_dump seq_loop_csv_dumper_220;
    seq_loop_monitor #(15) seq_loop_monitor_220;
    seq_loop_intf#(15) seq_loop_intf_221(clock,reset);
    assign seq_loop_intf_221.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state12;
    assign seq_loop_intf_221.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_221.pre_loop_state1 = 15'h0;
    assign seq_loop_intf_221.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_221.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state1;
    assign seq_loop_intf_221.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_221.post_loop_state1 = 15'h0;
    assign seq_loop_intf_221.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_221.post_loop_state2 = 15'h0;
    assign seq_loop_intf_221.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_221.post_loop_state3 = 15'h0;
    assign seq_loop_intf_221.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_221.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state14;
    assign seq_loop_intf_221.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_221.quit_loop_state1 = 15'h0;
    assign seq_loop_intf_221.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_221.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_CS_fsm;
    assign seq_loop_intf_221.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state14;
    assign seq_loop_intf_221.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_zint_bezout_1_fu_3626.grp_zint_co_reduce_mod_1_fu_674.ap_ST_fsm_state15;
    assign seq_loop_intf_221.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_221.iter_end_state1 = 15'h0;
    assign seq_loop_intf_221.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_221.one_state_loop = 1'b0;
    assign seq_loop_intf_221.one_state_block = 1'b0;
    assign seq_loop_intf_221.finish = finish;
    csv_file_dump seq_loop_csv_dumper_221;
    seq_loop_monitor #(15) seq_loop_monitor_221;
    seq_loop_intf#(7) seq_loop_intf_222(clock,reset);
    assign seq_loop_intf_222.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state5;
    assign seq_loop_intf_222.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_222.pre_loop_state1 = 7'h0;
    assign seq_loop_intf_222.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_222.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state4;
    assign seq_loop_intf_222.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_222.post_loop_state1 = 7'h0;
    assign seq_loop_intf_222.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_222.post_loop_state2 = 7'h0;
    assign seq_loop_intf_222.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_222.post_loop_state3 = 7'h0;
    assign seq_loop_intf_222.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_222.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state6;
    assign seq_loop_intf_222.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_222.quit_loop_state1 = 7'h0;
    assign seq_loop_intf_222.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_222.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_CS_fsm;
    assign seq_loop_intf_222.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state6;
    assign seq_loop_intf_222.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state7;
    assign seq_loop_intf_222.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_222.iter_end_state1 = 7'h0;
    assign seq_loop_intf_222.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_222.one_state_loop = 1'b0;
    assign seq_loop_intf_222.one_state_block = 1'b0;
    assign seq_loop_intf_222.finish = finish;
    csv_file_dump seq_loop_csv_dumper_222;
    seq_loop_monitor #(7) seq_loop_monitor_222;
    seq_loop_intf#(7) seq_loop_intf_223(clock,reset);
    assign seq_loop_intf_223.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state3;
    assign seq_loop_intf_223.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_223.pre_loop_state1 = 7'h0;
    assign seq_loop_intf_223.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_223.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state2;
    assign seq_loop_intf_223.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_223.post_loop_state1 = 7'h0;
    assign seq_loop_intf_223.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_223.post_loop_state2 = 7'h0;
    assign seq_loop_intf_223.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_223.post_loop_state3 = 7'h0;
    assign seq_loop_intf_223.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_223.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state4;
    assign seq_loop_intf_223.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_223.quit_loop_state1 = 7'h0;
    assign seq_loop_intf_223.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_223.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_CS_fsm;
    assign seq_loop_intf_223.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state4;
    assign seq_loop_intf_223.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state6;
    assign seq_loop_intf_223.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_223.iter_end_state1 = 7'h0;
    assign seq_loop_intf_223.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_223.one_state_loop = 1'b0;
    assign seq_loop_intf_223.one_state_block = 1'b0;
    assign seq_loop_intf_223.finish = finish;
    csv_file_dump seq_loop_csv_dumper_223;
    seq_loop_monitor #(7) seq_loop_monitor_223;
    seq_loop_intf#(7) seq_loop_intf_224(clock,reset);
    assign seq_loop_intf_224.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state1;
    assign seq_loop_intf_224.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_224.pre_loop_state1 = 7'h0;
    assign seq_loop_intf_224.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_224.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state1;
    assign seq_loop_intf_224.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_224.post_loop_state1 = 7'h0;
    assign seq_loop_intf_224.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_224.post_loop_state2 = 7'h0;
    assign seq_loop_intf_224.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_224.post_loop_state3 = 7'h0;
    assign seq_loop_intf_224.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_224.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state2;
    assign seq_loop_intf_224.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_224.quit_loop_state1 = 7'h0;
    assign seq_loop_intf_224.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_224.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_CS_fsm;
    assign seq_loop_intf_224.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state2;
    assign seq_loop_intf_224.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_1_fu_3632.ap_ST_fsm_state4;
    assign seq_loop_intf_224.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_224.iter_end_state1 = 7'h0;
    assign seq_loop_intf_224.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_224.one_state_loop = 1'b0;
    assign seq_loop_intf_224.one_state_block = 1'b0;
    assign seq_loop_intf_224.finish = finish;
    csv_file_dump seq_loop_csv_dumper_224;
    seq_loop_monitor #(7) seq_loop_monitor_224;
    seq_loop_intf#(44) seq_loop_intf_225(clock,reset);
    assign seq_loop_intf_225.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state8;
    assign seq_loop_intf_225.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_225.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_225.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_225.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state11;
    assign seq_loop_intf_225.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_225.post_loop_state1 = 44'h0;
    assign seq_loop_intf_225.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_225.post_loop_state2 = 44'h0;
    assign seq_loop_intf_225.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_225.post_loop_state3 = 44'h0;
    assign seq_loop_intf_225.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_225.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state9;
    assign seq_loop_intf_225.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_225.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_225.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_225.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_225.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state9;
    assign seq_loop_intf_225.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state10;
    assign seq_loop_intf_225.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_225.iter_end_state1 = 44'h0;
    assign seq_loop_intf_225.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_225.one_state_loop = 1'b0;
    assign seq_loop_intf_225.one_state_block = 1'b0;
    assign seq_loop_intf_225.finish = finish;
    csv_file_dump seq_loop_csv_dumper_225;
    seq_loop_monitor #(44) seq_loop_monitor_225;
    seq_loop_intf#(44) seq_loop_intf_226(clock,reset);
    assign seq_loop_intf_226.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state11;
    assign seq_loop_intf_226.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_226.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_226.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_226.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state13;
    assign seq_loop_intf_226.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_226.post_loop_state1 = 44'h0;
    assign seq_loop_intf_226.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_226.post_loop_state2 = 44'h0;
    assign seq_loop_intf_226.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_226.post_loop_state3 = 44'h0;
    assign seq_loop_intf_226.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_226.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state12;
    assign seq_loop_intf_226.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_226.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_226.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_226.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_226.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state12;
    assign seq_loop_intf_226.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state12;
    assign seq_loop_intf_226.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_226.iter_end_state1 = 44'h0;
    assign seq_loop_intf_226.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_226.one_state_loop = 1'b1;
    assign seq_loop_intf_226.one_state_block = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state12_blk;
    assign seq_loop_intf_226.finish = finish;
    csv_file_dump seq_loop_csv_dumper_226;
    seq_loop_monitor #(44) seq_loop_monitor_226;
    seq_loop_intf#(44) seq_loop_intf_227(clock,reset);
    assign seq_loop_intf_227.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state12;
    assign seq_loop_intf_227.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_227.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_227.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_227.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state15;
    assign seq_loop_intf_227.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_227.post_loop_state1 = 44'h0;
    assign seq_loop_intf_227.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_227.post_loop_state2 = 44'h0;
    assign seq_loop_intf_227.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_227.post_loop_state3 = 44'h0;
    assign seq_loop_intf_227.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_227.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state13;
    assign seq_loop_intf_227.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_227.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_227.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_227.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_227.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state13;
    assign seq_loop_intf_227.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state14;
    assign seq_loop_intf_227.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_227.iter_end_state1 = 44'h0;
    assign seq_loop_intf_227.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_227.one_state_loop = 1'b0;
    assign seq_loop_intf_227.one_state_block = 1'b0;
    assign seq_loop_intf_227.finish = finish;
    csv_file_dump seq_loop_csv_dumper_227;
    seq_loop_monitor #(44) seq_loop_monitor_227;
    seq_loop_intf#(44) seq_loop_intf_228(clock,reset);
    assign seq_loop_intf_228.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state15;
    assign seq_loop_intf_228.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_228.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_228.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_228.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state19;
    assign seq_loop_intf_228.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_228.post_loop_state1 = 44'h0;
    assign seq_loop_intf_228.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_228.post_loop_state2 = 44'h0;
    assign seq_loop_intf_228.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_228.post_loop_state3 = 44'h0;
    assign seq_loop_intf_228.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_228.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state16;
    assign seq_loop_intf_228.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_228.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_228.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_228.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_228.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state16;
    assign seq_loop_intf_228.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state18;
    assign seq_loop_intf_228.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_228.iter_end_state1 = 44'h0;
    assign seq_loop_intf_228.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_228.one_state_loop = 1'b0;
    assign seq_loop_intf_228.one_state_block = 1'b0;
    assign seq_loop_intf_228.finish = finish;
    csv_file_dump seq_loop_csv_dumper_228;
    seq_loop_monitor #(44) seq_loop_monitor_228;
    seq_loop_intf#(44) seq_loop_intf_229(clock,reset);
    assign seq_loop_intf_229.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state16;
    assign seq_loop_intf_229.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_229.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_229.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_229.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state21;
    assign seq_loop_intf_229.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_229.post_loop_state1 = 44'h0;
    assign seq_loop_intf_229.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_229.post_loop_state2 = 44'h0;
    assign seq_loop_intf_229.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_229.post_loop_state3 = 44'h0;
    assign seq_loop_intf_229.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_229.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state19;
    assign seq_loop_intf_229.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_229.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_229.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_229.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_229.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state19;
    assign seq_loop_intf_229.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state20;
    assign seq_loop_intf_229.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_229.iter_end_state1 = 44'h0;
    assign seq_loop_intf_229.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_229.one_state_loop = 1'b0;
    assign seq_loop_intf_229.one_state_block = 1'b0;
    assign seq_loop_intf_229.finish = finish;
    csv_file_dump seq_loop_csv_dumper_229;
    seq_loop_monitor #(44) seq_loop_monitor_229;
    seq_loop_intf#(44) seq_loop_intf_230(clock,reset);
    assign seq_loop_intf_230.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state22;
    assign seq_loop_intf_230.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_230.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_230.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_230.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state25;
    assign seq_loop_intf_230.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_230.post_loop_state1 = 44'h0;
    assign seq_loop_intf_230.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_230.post_loop_state2 = 44'h0;
    assign seq_loop_intf_230.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_230.post_loop_state3 = 44'h0;
    assign seq_loop_intf_230.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_230.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state24;
    assign seq_loop_intf_230.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_230.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_230.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_230.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_230.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state23;
    assign seq_loop_intf_230.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state24;
    assign seq_loop_intf_230.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_230.iter_end_state1 = 44'h0;
    assign seq_loop_intf_230.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_230.one_state_loop = 1'b0;
    assign seq_loop_intf_230.one_state_block = 1'b0;
    assign seq_loop_intf_230.finish = finish;
    csv_file_dump seq_loop_csv_dumper_230;
    seq_loop_monitor #(44) seq_loop_monitor_230;
    seq_loop_intf#(44) seq_loop_intf_231(clock,reset);
    assign seq_loop_intf_231.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state21;
    assign seq_loop_intf_231.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_231.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_231.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_231.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state26;
    assign seq_loop_intf_231.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_231.post_loop_state1 = 44'h0;
    assign seq_loop_intf_231.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_231.post_loop_state2 = 44'h0;
    assign seq_loop_intf_231.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_231.post_loop_state3 = 44'h0;
    assign seq_loop_intf_231.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_231.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state22;
    assign seq_loop_intf_231.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_231.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_231.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_231.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_231.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state22;
    assign seq_loop_intf_231.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state25;
    assign seq_loop_intf_231.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_231.iter_end_state1 = 44'h0;
    assign seq_loop_intf_231.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_231.one_state_loop = 1'b0;
    assign seq_loop_intf_231.one_state_block = 1'b0;
    assign seq_loop_intf_231.finish = finish;
    csv_file_dump seq_loop_csv_dumper_231;
    seq_loop_monitor #(44) seq_loop_monitor_231;
    seq_loop_intf#(44) seq_loop_intf_232(clock,reset);
    assign seq_loop_intf_232.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state26;
    assign seq_loop_intf_232.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_232.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_232.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_232.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state30;
    assign seq_loop_intf_232.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_232.post_loop_state1 = 44'h0;
    assign seq_loop_intf_232.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_232.post_loop_state2 = 44'h0;
    assign seq_loop_intf_232.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_232.post_loop_state3 = 44'h0;
    assign seq_loop_intf_232.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_232.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state27;
    assign seq_loop_intf_232.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_232.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_232.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_232.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_232.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state27;
    assign seq_loop_intf_232.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state29;
    assign seq_loop_intf_232.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_232.iter_end_state1 = 44'h0;
    assign seq_loop_intf_232.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_232.one_state_loop = 1'b0;
    assign seq_loop_intf_232.one_state_block = 1'b0;
    assign seq_loop_intf_232.finish = finish;
    csv_file_dump seq_loop_csv_dumper_232;
    seq_loop_monitor #(44) seq_loop_monitor_232;
    seq_loop_intf#(44) seq_loop_intf_233(clock,reset);
    assign seq_loop_intf_233.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state34;
    assign seq_loop_intf_233.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_233.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_233.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_233.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state31;
    assign seq_loop_intf_233.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_233.post_loop_state1 = 44'h0;
    assign seq_loop_intf_233.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_233.post_loop_state2 = 44'h0;
    assign seq_loop_intf_233.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_233.post_loop_state3 = 44'h0;
    assign seq_loop_intf_233.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_233.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state35;
    assign seq_loop_intf_233.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_233.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_233.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_233.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_233.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state35;
    assign seq_loop_intf_233.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state37;
    assign seq_loop_intf_233.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_233.iter_end_state1 = 44'h0;
    assign seq_loop_intf_233.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_233.one_state_loop = 1'b0;
    assign seq_loop_intf_233.one_state_block = 1'b0;
    assign seq_loop_intf_233.finish = finish;
    csv_file_dump seq_loop_csv_dumper_233;
    seq_loop_monitor #(44) seq_loop_monitor_233;
    seq_loop_intf#(44) seq_loop_intf_234(clock,reset);
    assign seq_loop_intf_234.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state30;
    assign seq_loop_intf_234.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_234.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_234.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_234.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state30;
    assign seq_loop_intf_234.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_234.post_loop_state1 = 44'h0;
    assign seq_loop_intf_234.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_234.post_loop_state2 = 44'h0;
    assign seq_loop_intf_234.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_234.post_loop_state3 = 44'h0;
    assign seq_loop_intf_234.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_234.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state31;
    assign seq_loop_intf_234.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_234.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_234.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_234.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_234.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state31;
    assign seq_loop_intf_234.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state35;
    assign seq_loop_intf_234.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_234.iter_end_state1 = 44'h0;
    assign seq_loop_intf_234.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_234.one_state_loop = 1'b0;
    assign seq_loop_intf_234.one_state_block = 1'b0;
    assign seq_loop_intf_234.finish = finish;
    csv_file_dump seq_loop_csv_dumper_234;
    seq_loop_monitor #(44) seq_loop_monitor_234;
    seq_loop_intf#(44) seq_loop_intf_235(clock,reset);
    assign seq_loop_intf_235.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state27;
    assign seq_loop_intf_235.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_235.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_235.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_235.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state38;
    assign seq_loop_intf_235.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_235.post_loop_state1 = 44'h0;
    assign seq_loop_intf_235.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_235.post_loop_state2 = 44'h0;
    assign seq_loop_intf_235.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_235.post_loop_state3 = 44'h0;
    assign seq_loop_intf_235.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_235.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state30;
    assign seq_loop_intf_235.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_235.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_235.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_235.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_235.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state30;
    assign seq_loop_intf_235.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state31;
    assign seq_loop_intf_235.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_235.iter_end_state1 = 44'h0;
    assign seq_loop_intf_235.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_235.one_state_loop = 1'b0;
    assign seq_loop_intf_235.one_state_block = 1'b0;
    assign seq_loop_intf_235.finish = finish;
    csv_file_dump seq_loop_csv_dumper_235;
    seq_loop_monitor #(44) seq_loop_monitor_235;
    seq_loop_intf#(44) seq_loop_intf_236(clock,reset);
    assign seq_loop_intf_236.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state30;
    assign seq_loop_intf_236.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_236.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_236.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_236.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state2;
    assign seq_loop_intf_236.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_236.post_loop_state1 = 44'h0;
    assign seq_loop_intf_236.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_236.post_loop_state2 = 44'h0;
    assign seq_loop_intf_236.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_236.post_loop_state3 = 44'h0;
    assign seq_loop_intf_236.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_236.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state38;
    assign seq_loop_intf_236.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_236.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_236.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_236.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_236.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state38;
    assign seq_loop_intf_236.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state39;
    assign seq_loop_intf_236.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_236.iter_end_state1 = 44'h0;
    assign seq_loop_intf_236.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_236.one_state_loop = 1'b0;
    assign seq_loop_intf_236.one_state_block = 1'b0;
    assign seq_loop_intf_236.finish = finish;
    csv_file_dump seq_loop_csv_dumper_236;
    seq_loop_monitor #(44) seq_loop_monitor_236;
    seq_loop_intf#(44) seq_loop_intf_237(clock,reset);
    assign seq_loop_intf_237.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state1;
    assign seq_loop_intf_237.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_237.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_237.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_237.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state40;
    assign seq_loop_intf_237.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_237.post_loop_state1 = 44'h0;
    assign seq_loop_intf_237.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_237.post_loop_state2 = 44'h0;
    assign seq_loop_intf_237.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_237.post_loop_state3 = 44'h0;
    assign seq_loop_intf_237.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_237.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state2;
    assign seq_loop_intf_237.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_237.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_237.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_237.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_237.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state2;
    assign seq_loop_intf_237.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state38;
    assign seq_loop_intf_237.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_237.iter_end_state1 = 44'h0;
    assign seq_loop_intf_237.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_237.one_state_loop = 1'b0;
    assign seq_loop_intf_237.one_state_block = 1'b0;
    assign seq_loop_intf_237.finish = finish;
    csv_file_dump seq_loop_csv_dumper_237;
    seq_loop_monitor #(44) seq_loop_monitor_237;
    seq_loop_intf#(44) seq_loop_intf_238(clock,reset);
    assign seq_loop_intf_238.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state42;
    assign seq_loop_intf_238.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_238.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_238.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_238.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state41;
    assign seq_loop_intf_238.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_238.post_loop_state1 = 44'h0;
    assign seq_loop_intf_238.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_238.post_loop_state2 = 44'h0;
    assign seq_loop_intf_238.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_238.post_loop_state3 = 44'h0;
    assign seq_loop_intf_238.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_238.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state43;
    assign seq_loop_intf_238.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_238.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_238.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_238.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_238.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state43;
    assign seq_loop_intf_238.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state44;
    assign seq_loop_intf_238.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_238.iter_end_state1 = 44'h0;
    assign seq_loop_intf_238.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_238.one_state_loop = 1'b0;
    assign seq_loop_intf_238.one_state_block = 1'b0;
    assign seq_loop_intf_238.finish = finish;
    csv_file_dump seq_loop_csv_dumper_238;
    seq_loop_monitor #(44) seq_loop_monitor_238;
    seq_loop_intf#(44) seq_loop_intf_239(clock,reset);
    assign seq_loop_intf_239.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state40;
    assign seq_loop_intf_239.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_239.pre_loop_state1 = 44'h0;
    assign seq_loop_intf_239.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_239.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state1;
    assign seq_loop_intf_239.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_239.post_loop_state1 = 44'h0;
    assign seq_loop_intf_239.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_239.post_loop_state2 = 44'h0;
    assign seq_loop_intf_239.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_239.post_loop_state3 = 44'h0;
    assign seq_loop_intf_239.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_239.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state41;
    assign seq_loop_intf_239.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_239.quit_loop_state1 = 44'h0;
    assign seq_loop_intf_239.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_239.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_CS_fsm;
    assign seq_loop_intf_239.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state41;
    assign seq_loop_intf_239.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.ap_ST_fsm_state43;
    assign seq_loop_intf_239.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_239.iter_end_state1 = 44'h0;
    assign seq_loop_intf_239.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_239.one_state_loop = 1'b0;
    assign seq_loop_intf_239.one_state_block = 1'b0;
    assign seq_loop_intf_239.finish = finish;
    csv_file_dump seq_loop_csv_dumper_239;
    seq_loop_monitor #(44) seq_loop_monitor_239;
    seq_loop_intf#(19) seq_loop_intf_240(clock,reset);
    assign seq_loop_intf_240.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state8;
    assign seq_loop_intf_240.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_240.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_240.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_240.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state11;
    assign seq_loop_intf_240.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_240.post_loop_state1 = 19'h0;
    assign seq_loop_intf_240.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_240.post_loop_state2 = 19'h0;
    assign seq_loop_intf_240.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_240.post_loop_state3 = 19'h0;
    assign seq_loop_intf_240.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_240.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state10;
    assign seq_loop_intf_240.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_240.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_240.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_240.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_CS_fsm;
    assign seq_loop_intf_240.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state9;
    assign seq_loop_intf_240.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state10;
    assign seq_loop_intf_240.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_240.iter_end_state1 = 19'h0;
    assign seq_loop_intf_240.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_240.one_state_loop = 1'b0;
    assign seq_loop_intf_240.one_state_block = 1'b0;
    assign seq_loop_intf_240.finish = finish;
    csv_file_dump seq_loop_csv_dumper_240;
    seq_loop_monitor #(19) seq_loop_monitor_240;
    seq_loop_intf#(19) seq_loop_intf_241(clock,reset);
    assign seq_loop_intf_241.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state10;
    assign seq_loop_intf_241.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_241.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_241.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_241.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state7;
    assign seq_loop_intf_241.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_241.post_loop_state1 = 19'h0;
    assign seq_loop_intf_241.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_241.post_loop_state2 = 19'h0;
    assign seq_loop_intf_241.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_241.post_loop_state3 = 19'h0;
    assign seq_loop_intf_241.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_241.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state11;
    assign seq_loop_intf_241.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_241.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_241.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_241.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_CS_fsm;
    assign seq_loop_intf_241.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state11;
    assign seq_loop_intf_241.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state12;
    assign seq_loop_intf_241.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_241.iter_end_state1 = 19'h0;
    assign seq_loop_intf_241.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_241.one_state_loop = 1'b0;
    assign seq_loop_intf_241.one_state_block = 1'b0;
    assign seq_loop_intf_241.finish = finish;
    csv_file_dump seq_loop_csv_dumper_241;
    seq_loop_monitor #(19) seq_loop_monitor_241;
    seq_loop_intf#(19) seq_loop_intf_242(clock,reset);
    assign seq_loop_intf_242.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state6;
    assign seq_loop_intf_242.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_242.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_242.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_242.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state13;
    assign seq_loop_intf_242.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_242.post_loop_state1 = 19'h0;
    assign seq_loop_intf_242.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_242.post_loop_state2 = 19'h0;
    assign seq_loop_intf_242.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_242.post_loop_state3 = 19'h0;
    assign seq_loop_intf_242.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_242.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state7;
    assign seq_loop_intf_242.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_242.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_242.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_242.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_CS_fsm;
    assign seq_loop_intf_242.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state7;
    assign seq_loop_intf_242.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state11;
    assign seq_loop_intf_242.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_242.iter_end_state1 = 19'h0;
    assign seq_loop_intf_242.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_242.one_state_loop = 1'b0;
    assign seq_loop_intf_242.one_state_block = 1'b0;
    assign seq_loop_intf_242.finish = finish;
    csv_file_dump seq_loop_csv_dumper_242;
    seq_loop_monitor #(19) seq_loop_monitor_242;
    seq_loop_intf#(19) seq_loop_intf_243(clock,reset);
    assign seq_loop_intf_243.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state7;
    assign seq_loop_intf_243.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_243.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_243.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_243.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state2;
    assign seq_loop_intf_243.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_243.post_loop_state1 = 19'h0;
    assign seq_loop_intf_243.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_243.post_loop_state2 = 19'h0;
    assign seq_loop_intf_243.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_243.post_loop_state3 = 19'h0;
    assign seq_loop_intf_243.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_243.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state13;
    assign seq_loop_intf_243.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_243.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_243.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_243.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_CS_fsm;
    assign seq_loop_intf_243.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state13;
    assign seq_loop_intf_243.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state14;
    assign seq_loop_intf_243.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_243.iter_end_state1 = 19'h0;
    assign seq_loop_intf_243.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_243.one_state_loop = 1'b0;
    assign seq_loop_intf_243.one_state_block = 1'b0;
    assign seq_loop_intf_243.finish = finish;
    csv_file_dump seq_loop_csv_dumper_243;
    seq_loop_monitor #(19) seq_loop_monitor_243;
    seq_loop_intf#(19) seq_loop_intf_244(clock,reset);
    assign seq_loop_intf_244.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state1;
    assign seq_loop_intf_244.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_244.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_244.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_244.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state15;
    assign seq_loop_intf_244.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_244.post_loop_state1 = 19'h0;
    assign seq_loop_intf_244.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_244.post_loop_state2 = 19'h0;
    assign seq_loop_intf_244.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_244.post_loop_state3 = 19'h0;
    assign seq_loop_intf_244.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_244.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state2;
    assign seq_loop_intf_244.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_244.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_244.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_244.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_CS_fsm;
    assign seq_loop_intf_244.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state2;
    assign seq_loop_intf_244.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state13;
    assign seq_loop_intf_244.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_244.iter_end_state1 = 19'h0;
    assign seq_loop_intf_244.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_244.one_state_loop = 1'b0;
    assign seq_loop_intf_244.one_state_block = 1'b0;
    assign seq_loop_intf_244.finish = finish;
    csv_file_dump seq_loop_csv_dumper_244;
    seq_loop_monitor #(19) seq_loop_monitor_244;
    seq_loop_intf#(19) seq_loop_intf_245(clock,reset);
    assign seq_loop_intf_245.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state15;
    assign seq_loop_intf_245.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_245.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_245.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_245.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state18;
    assign seq_loop_intf_245.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_245.post_loop_state1 = 19'h0;
    assign seq_loop_intf_245.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_245.post_loop_state2 = 19'h0;
    assign seq_loop_intf_245.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_245.post_loop_state3 = 19'h0;
    assign seq_loop_intf_245.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_245.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state17;
    assign seq_loop_intf_245.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_245.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_245.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_245.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_CS_fsm;
    assign seq_loop_intf_245.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state16;
    assign seq_loop_intf_245.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state17;
    assign seq_loop_intf_245.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_245.iter_end_state1 = 19'h0;
    assign seq_loop_intf_245.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_245.one_state_loop = 1'b0;
    assign seq_loop_intf_245.one_state_block = 1'b0;
    assign seq_loop_intf_245.finish = finish;
    csv_file_dump seq_loop_csv_dumper_245;
    seq_loop_monitor #(19) seq_loop_monitor_245;
    seq_loop_intf#(19) seq_loop_intf_246(clock,reset);
    assign seq_loop_intf_246.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state17;
    assign seq_loop_intf_246.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_246.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_246.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_246.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state15;
    assign seq_loop_intf_246.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_246.post_loop_state1 = 19'h0;
    assign seq_loop_intf_246.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_246.post_loop_state2 = 19'h0;
    assign seq_loop_intf_246.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_246.post_loop_state3 = 19'h0;
    assign seq_loop_intf_246.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_246.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state18;
    assign seq_loop_intf_246.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_246.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_246.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_246.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_CS_fsm;
    assign seq_loop_intf_246.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state18;
    assign seq_loop_intf_246.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state19;
    assign seq_loop_intf_246.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_246.iter_end_state1 = 19'h0;
    assign seq_loop_intf_246.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_246.one_state_loop = 1'b0;
    assign seq_loop_intf_246.one_state_block = 1'b0;
    assign seq_loop_intf_246.finish = finish;
    csv_file_dump seq_loop_csv_dumper_246;
    seq_loop_monitor #(19) seq_loop_monitor_246;
    seq_loop_intf#(19) seq_loop_intf_247(clock,reset);
    assign seq_loop_intf_247.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state2;
    assign seq_loop_intf_247.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_247.pre_loop_state1 = 19'h0;
    assign seq_loop_intf_247.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_247.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state1;
    assign seq_loop_intf_247.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_247.post_loop_state1 = 19'h0;
    assign seq_loop_intf_247.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_247.post_loop_state2 = 19'h0;
    assign seq_loop_intf_247.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_247.post_loop_state3 = 19'h0;
    assign seq_loop_intf_247.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_247.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state15;
    assign seq_loop_intf_247.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_247.quit_loop_state1 = 19'h0;
    assign seq_loop_intf_247.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_247.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_CS_fsm;
    assign seq_loop_intf_247.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state15;
    assign seq_loop_intf_247.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_zint_rebuild_CRT_1_fu_1154.ap_ST_fsm_state18;
    assign seq_loop_intf_247.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_247.iter_end_state1 = 19'h0;
    assign seq_loop_intf_247.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_247.one_state_loop = 1'b0;
    assign seq_loop_intf_247.one_state_block = 1'b0;
    assign seq_loop_intf_247.finish = finish;
    csv_file_dump seq_loop_csv_dumper_247;
    seq_loop_monitor #(19) seq_loop_monitor_247;
    seq_loop_intf#(9) seq_loop_intf_248(clock,reset);
    assign seq_loop_intf_248.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state6;
    assign seq_loop_intf_248.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_248.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_248.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_248.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state3;
    assign seq_loop_intf_248.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_248.post_loop_state1 = 9'h0;
    assign seq_loop_intf_248.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_248.post_loop_state2 = 9'h0;
    assign seq_loop_intf_248.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_248.post_loop_state3 = 9'h0;
    assign seq_loop_intf_248.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_248.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state7;
    assign seq_loop_intf_248.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_248.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_248.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_248.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_CS_fsm;
    assign seq_loop_intf_248.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state7;
    assign seq_loop_intf_248.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state9;
    assign seq_loop_intf_248.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_248.iter_end_state1 = 9'h0;
    assign seq_loop_intf_248.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_248.one_state_loop = 1'b0;
    assign seq_loop_intf_248.one_state_block = 1'b0;
    assign seq_loop_intf_248.finish = finish;
    csv_file_dump seq_loop_csv_dumper_248;
    seq_loop_monitor #(9) seq_loop_monitor_248;
    seq_loop_intf#(9) seq_loop_intf_249(clock,reset);
    assign seq_loop_intf_249.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state2;
    assign seq_loop_intf_249.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_249.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_249.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_249.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state2;
    assign seq_loop_intf_249.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_249.post_loop_state1 = 9'h0;
    assign seq_loop_intf_249.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_249.post_loop_state2 = 9'h0;
    assign seq_loop_intf_249.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_249.post_loop_state3 = 9'h0;
    assign seq_loop_intf_249.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_249.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state3;
    assign seq_loop_intf_249.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_249.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_249.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_249.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_CS_fsm;
    assign seq_loop_intf_249.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state3;
    assign seq_loop_intf_249.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state7;
    assign seq_loop_intf_249.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_249.iter_end_state1 = 9'h0;
    assign seq_loop_intf_249.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_249.one_state_loop = 1'b0;
    assign seq_loop_intf_249.one_state_block = 1'b0;
    assign seq_loop_intf_249.finish = finish;
    csv_file_dump seq_loop_csv_dumper_249;
    seq_loop_monitor #(9) seq_loop_monitor_249;
    seq_loop_intf#(9) seq_loop_intf_250(clock,reset);
    assign seq_loop_intf_250.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state1;
    assign seq_loop_intf_250.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_250.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_250.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_250.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state1;
    assign seq_loop_intf_250.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_250.post_loop_state1 = 9'h0;
    assign seq_loop_intf_250.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_250.post_loop_state2 = 9'h0;
    assign seq_loop_intf_250.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_250.post_loop_state3 = 9'h0;
    assign seq_loop_intf_250.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_250.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state2;
    assign seq_loop_intf_250.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_250.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_250.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_250.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_CS_fsm;
    assign seq_loop_intf_250.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state2;
    assign seq_loop_intf_250.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_solve_NTRU_all_1_fu_478.grp_poly_sub_scaled_ntt_1_fu_3649.grp_modp_NTT2_ext_1_fu_1171.ap_ST_fsm_state3;
    assign seq_loop_intf_250.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_250.iter_end_state1 = 9'h0;
    assign seq_loop_intf_250.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_250.one_state_loop = 1'b0;
    assign seq_loop_intf_250.one_state_block = 1'b0;
    assign seq_loop_intf_250.finish = finish;
    csv_file_dump seq_loop_csv_dumper_250;
    seq_loop_monitor #(9) seq_loop_monitor_250;
    seq_loop_intf#(9) seq_loop_intf_251(clock,reset);
    assign seq_loop_intf_251.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state6;
    assign seq_loop_intf_251.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_251.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_251.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_251.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state3;
    assign seq_loop_intf_251.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_251.post_loop_state1 = 9'h0;
    assign seq_loop_intf_251.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_251.post_loop_state2 = 9'h0;
    assign seq_loop_intf_251.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_251.post_loop_state3 = 9'h0;
    assign seq_loop_intf_251.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_251.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state7;
    assign seq_loop_intf_251.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_251.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_251.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_251.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_CS_fsm;
    assign seq_loop_intf_251.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state7;
    assign seq_loop_intf_251.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state9;
    assign seq_loop_intf_251.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_251.iter_end_state1 = 9'h0;
    assign seq_loop_intf_251.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_251.one_state_loop = 1'b0;
    assign seq_loop_intf_251.one_state_block = 1'b0;
    assign seq_loop_intf_251.finish = finish;
    csv_file_dump seq_loop_csv_dumper_251;
    seq_loop_monitor #(9) seq_loop_monitor_251;
    seq_loop_intf#(9) seq_loop_intf_252(clock,reset);
    assign seq_loop_intf_252.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state2;
    assign seq_loop_intf_252.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_252.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_252.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_252.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state2;
    assign seq_loop_intf_252.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_252.post_loop_state1 = 9'h0;
    assign seq_loop_intf_252.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_252.post_loop_state2 = 9'h0;
    assign seq_loop_intf_252.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_252.post_loop_state3 = 9'h0;
    assign seq_loop_intf_252.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_252.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state3;
    assign seq_loop_intf_252.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_252.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_252.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_252.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_CS_fsm;
    assign seq_loop_intf_252.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state3;
    assign seq_loop_intf_252.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state7;
    assign seq_loop_intf_252.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_252.iter_end_state1 = 9'h0;
    assign seq_loop_intf_252.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_252.one_state_loop = 1'b0;
    assign seq_loop_intf_252.one_state_block = 1'b0;
    assign seq_loop_intf_252.finish = finish;
    csv_file_dump seq_loop_csv_dumper_252;
    seq_loop_monitor #(9) seq_loop_monitor_252;
    seq_loop_intf#(9) seq_loop_intf_253(clock,reset);
    assign seq_loop_intf_253.pre_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state1;
    assign seq_loop_intf_253.pre_states_valid[0] = 1'b1;
    assign seq_loop_intf_253.pre_loop_state1 = 9'h0;
    assign seq_loop_intf_253.pre_states_valid[1] = 1'b0;
    assign seq_loop_intf_253.post_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state1;
    assign seq_loop_intf_253.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_253.post_loop_state1 = 9'h0;
    assign seq_loop_intf_253.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_253.post_loop_state2 = 9'h0;
    assign seq_loop_intf_253.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_253.post_loop_state3 = 9'h0;
    assign seq_loop_intf_253.post_states_valid[3] = 1'b0;
    assign seq_loop_intf_253.quit_loop_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state2;
    assign seq_loop_intf_253.quit_states_valid[0] = 1'b1;
    assign seq_loop_intf_253.quit_loop_state1 = 9'h0;
    assign seq_loop_intf_253.quit_states_valid[1] = 1'b0;
    assign seq_loop_intf_253.cur_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_CS_fsm;
    assign seq_loop_intf_253.iter_start_state = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state2;
    assign seq_loop_intf_253.iter_end_state0 = AESL_inst_keygen.grp_solve_NTRU_fu_1364.grp_modp_NTT2_ext_1_fu_542.ap_ST_fsm_state3;
    assign seq_loop_intf_253.iter_end_states_valid[0] = 1'b1;
    assign seq_loop_intf_253.iter_end_state1 = 9'h0;
    assign seq_loop_intf_253.iter_end_states_valid[1] = 1'b0;
    assign seq_loop_intf_253.one_state_loop = 1'b0;
    assign seq_loop_intf_253.one_state_block = 1'b0;
    assign seq_loop_intf_253.finish = finish;
    csv_file_dump seq_loop_csv_dumper_253;
    seq_loop_monitor #(9) seq_loop_monitor_253;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);
    mstatus_csv_dumper_7 = new("./module_status7.csv");
    module_monitor_7 = new(module_intf_7,mstatus_csv_dumper_7);
    mstatus_csv_dumper_8 = new("./module_status8.csv");
    module_monitor_8 = new(module_intf_8,mstatus_csv_dumper_8);
    mstatus_csv_dumper_9 = new("./module_status9.csv");
    module_monitor_9 = new(module_intf_9,mstatus_csv_dumper_9);
    mstatus_csv_dumper_10 = new("./module_status10.csv");
    module_monitor_10 = new(module_intf_10,mstatus_csv_dumper_10);
    mstatus_csv_dumper_11 = new("./module_status11.csv");
    module_monitor_11 = new(module_intf_11,mstatus_csv_dumper_11);
    mstatus_csv_dumper_12 = new("./module_status12.csv");
    module_monitor_12 = new(module_intf_12,mstatus_csv_dumper_12);
    mstatus_csv_dumper_13 = new("./module_status13.csv");
    module_monitor_13 = new(module_intf_13,mstatus_csv_dumper_13);
    mstatus_csv_dumper_14 = new("./module_status14.csv");
    module_monitor_14 = new(module_intf_14,mstatus_csv_dumper_14);
    mstatus_csv_dumper_15 = new("./module_status15.csv");
    module_monitor_15 = new(module_intf_15,mstatus_csv_dumper_15);
    mstatus_csv_dumper_16 = new("./module_status16.csv");
    module_monitor_16 = new(module_intf_16,mstatus_csv_dumper_16);
    mstatus_csv_dumper_17 = new("./module_status17.csv");
    module_monitor_17 = new(module_intf_17,mstatus_csv_dumper_17);
    mstatus_csv_dumper_18 = new("./module_status18.csv");
    module_monitor_18 = new(module_intf_18,mstatus_csv_dumper_18);
    mstatus_csv_dumper_19 = new("./module_status19.csv");
    module_monitor_19 = new(module_intf_19,mstatus_csv_dumper_19);
    mstatus_csv_dumper_20 = new("./module_status20.csv");
    module_monitor_20 = new(module_intf_20,mstatus_csv_dumper_20);
    mstatus_csv_dumper_21 = new("./module_status21.csv");
    module_monitor_21 = new(module_intf_21,mstatus_csv_dumper_21);
    mstatus_csv_dumper_22 = new("./module_status22.csv");
    module_monitor_22 = new(module_intf_22,mstatus_csv_dumper_22);
    mstatus_csv_dumper_23 = new("./module_status23.csv");
    module_monitor_23 = new(module_intf_23,mstatus_csv_dumper_23);
    mstatus_csv_dumper_24 = new("./module_status24.csv");
    module_monitor_24 = new(module_intf_24,mstatus_csv_dumper_24);
    mstatus_csv_dumper_25 = new("./module_status25.csv");
    module_monitor_25 = new(module_intf_25,mstatus_csv_dumper_25);
    mstatus_csv_dumper_26 = new("./module_status26.csv");
    module_monitor_26 = new(module_intf_26,mstatus_csv_dumper_26);
    mstatus_csv_dumper_27 = new("./module_status27.csv");
    module_monitor_27 = new(module_intf_27,mstatus_csv_dumper_27);
    mstatus_csv_dumper_28 = new("./module_status28.csv");
    module_monitor_28 = new(module_intf_28,mstatus_csv_dumper_28);
    mstatus_csv_dumper_29 = new("./module_status29.csv");
    module_monitor_29 = new(module_intf_29,mstatus_csv_dumper_29);
    mstatus_csv_dumper_30 = new("./module_status30.csv");
    module_monitor_30 = new(module_intf_30,mstatus_csv_dumper_30);
    mstatus_csv_dumper_31 = new("./module_status31.csv");
    module_monitor_31 = new(module_intf_31,mstatus_csv_dumper_31);
    mstatus_csv_dumper_32 = new("./module_status32.csv");
    module_monitor_32 = new(module_intf_32,mstatus_csv_dumper_32);
    mstatus_csv_dumper_33 = new("./module_status33.csv");
    module_monitor_33 = new(module_intf_33,mstatus_csv_dumper_33);
    mstatus_csv_dumper_34 = new("./module_status34.csv");
    module_monitor_34 = new(module_intf_34,mstatus_csv_dumper_34);
    mstatus_csv_dumper_35 = new("./module_status35.csv");
    module_monitor_35 = new(module_intf_35,mstatus_csv_dumper_35);
    mstatus_csv_dumper_36 = new("./module_status36.csv");
    module_monitor_36 = new(module_intf_36,mstatus_csv_dumper_36);
    mstatus_csv_dumper_37 = new("./module_status37.csv");
    module_monitor_37 = new(module_intf_37,mstatus_csv_dumper_37);
    mstatus_csv_dumper_38 = new("./module_status38.csv");
    module_monitor_38 = new(module_intf_38,mstatus_csv_dumper_38);
    mstatus_csv_dumper_39 = new("./module_status39.csv");
    module_monitor_39 = new(module_intf_39,mstatus_csv_dumper_39);
    mstatus_csv_dumper_40 = new("./module_status40.csv");
    module_monitor_40 = new(module_intf_40,mstatus_csv_dumper_40);
    mstatus_csv_dumper_41 = new("./module_status41.csv");
    module_monitor_41 = new(module_intf_41,mstatus_csv_dumper_41);
    mstatus_csv_dumper_42 = new("./module_status42.csv");
    module_monitor_42 = new(module_intf_42,mstatus_csv_dumper_42);
    mstatus_csv_dumper_43 = new("./module_status43.csv");
    module_monitor_43 = new(module_intf_43,mstatus_csv_dumper_43);
    mstatus_csv_dumper_44 = new("./module_status44.csv");
    module_monitor_44 = new(module_intf_44,mstatus_csv_dumper_44);
    mstatus_csv_dumper_45 = new("./module_status45.csv");
    module_monitor_45 = new(module_intf_45,mstatus_csv_dumper_45);
    mstatus_csv_dumper_46 = new("./module_status46.csv");
    module_monitor_46 = new(module_intf_46,mstatus_csv_dumper_46);
    mstatus_csv_dumper_47 = new("./module_status47.csv");
    module_monitor_47 = new(module_intf_47,mstatus_csv_dumper_47);
    mstatus_csv_dumper_48 = new("./module_status48.csv");
    module_monitor_48 = new(module_intf_48,mstatus_csv_dumper_48);
    mstatus_csv_dumper_49 = new("./module_status49.csv");
    module_monitor_49 = new(module_intf_49,mstatus_csv_dumper_49);
    mstatus_csv_dumper_50 = new("./module_status50.csv");
    module_monitor_50 = new(module_intf_50,mstatus_csv_dumper_50);
    mstatus_csv_dumper_51 = new("./module_status51.csv");
    module_monitor_51 = new(module_intf_51,mstatus_csv_dumper_51);
    mstatus_csv_dumper_52 = new("./module_status52.csv");
    module_monitor_52 = new(module_intf_52,mstatus_csv_dumper_52);
    mstatus_csv_dumper_53 = new("./module_status53.csv");
    module_monitor_53 = new(module_intf_53,mstatus_csv_dumper_53);
    mstatus_csv_dumper_54 = new("./module_status54.csv");
    module_monitor_54 = new(module_intf_54,mstatus_csv_dumper_54);
    mstatus_csv_dumper_55 = new("./module_status55.csv");
    module_monitor_55 = new(module_intf_55,mstatus_csv_dumper_55);
    mstatus_csv_dumper_56 = new("./module_status56.csv");
    module_monitor_56 = new(module_intf_56,mstatus_csv_dumper_56);
    mstatus_csv_dumper_57 = new("./module_status57.csv");
    module_monitor_57 = new(module_intf_57,mstatus_csv_dumper_57);
    mstatus_csv_dumper_58 = new("./module_status58.csv");
    module_monitor_58 = new(module_intf_58,mstatus_csv_dumper_58);
    mstatus_csv_dumper_59 = new("./module_status59.csv");
    module_monitor_59 = new(module_intf_59,mstatus_csv_dumper_59);
    mstatus_csv_dumper_60 = new("./module_status60.csv");
    module_monitor_60 = new(module_intf_60,mstatus_csv_dumper_60);
    mstatus_csv_dumper_61 = new("./module_status61.csv");
    module_monitor_61 = new(module_intf_61,mstatus_csv_dumper_61);
    mstatus_csv_dumper_62 = new("./module_status62.csv");
    module_monitor_62 = new(module_intf_62,mstatus_csv_dumper_62);
    mstatus_csv_dumper_63 = new("./module_status63.csv");
    module_monitor_63 = new(module_intf_63,mstatus_csv_dumper_63);
    mstatus_csv_dumper_64 = new("./module_status64.csv");
    module_monitor_64 = new(module_intf_64,mstatus_csv_dumper_64);
    mstatus_csv_dumper_65 = new("./module_status65.csv");
    module_monitor_65 = new(module_intf_65,mstatus_csv_dumper_65);
    mstatus_csv_dumper_66 = new("./module_status66.csv");
    module_monitor_66 = new(module_intf_66,mstatus_csv_dumper_66);
    mstatus_csv_dumper_67 = new("./module_status67.csv");
    module_monitor_67 = new(module_intf_67,mstatus_csv_dumper_67);



    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);
    seq_loop_csv_dumper_7 = new("./seq_loop_status7.csv");
    seq_loop_monitor_7 = new(seq_loop_intf_7,seq_loop_csv_dumper_7);
    seq_loop_csv_dumper_8 = new("./seq_loop_status8.csv");
    seq_loop_monitor_8 = new(seq_loop_intf_8,seq_loop_csv_dumper_8);
    seq_loop_csv_dumper_9 = new("./seq_loop_status9.csv");
    seq_loop_monitor_9 = new(seq_loop_intf_9,seq_loop_csv_dumper_9);
    seq_loop_csv_dumper_10 = new("./seq_loop_status10.csv");
    seq_loop_monitor_10 = new(seq_loop_intf_10,seq_loop_csv_dumper_10);
    seq_loop_csv_dumper_11 = new("./seq_loop_status11.csv");
    seq_loop_monitor_11 = new(seq_loop_intf_11,seq_loop_csv_dumper_11);
    seq_loop_csv_dumper_12 = new("./seq_loop_status12.csv");
    seq_loop_monitor_12 = new(seq_loop_intf_12,seq_loop_csv_dumper_12);
    seq_loop_csv_dumper_13 = new("./seq_loop_status13.csv");
    seq_loop_monitor_13 = new(seq_loop_intf_13,seq_loop_csv_dumper_13);
    seq_loop_csv_dumper_14 = new("./seq_loop_status14.csv");
    seq_loop_monitor_14 = new(seq_loop_intf_14,seq_loop_csv_dumper_14);
    seq_loop_csv_dumper_15 = new("./seq_loop_status15.csv");
    seq_loop_monitor_15 = new(seq_loop_intf_15,seq_loop_csv_dumper_15);
    seq_loop_csv_dumper_16 = new("./seq_loop_status16.csv");
    seq_loop_monitor_16 = new(seq_loop_intf_16,seq_loop_csv_dumper_16);
    seq_loop_csv_dumper_17 = new("./seq_loop_status17.csv");
    seq_loop_monitor_17 = new(seq_loop_intf_17,seq_loop_csv_dumper_17);
    seq_loop_csv_dumper_18 = new("./seq_loop_status18.csv");
    seq_loop_monitor_18 = new(seq_loop_intf_18,seq_loop_csv_dumper_18);
    seq_loop_csv_dumper_19 = new("./seq_loop_status19.csv");
    seq_loop_monitor_19 = new(seq_loop_intf_19,seq_loop_csv_dumper_19);
    seq_loop_csv_dumper_20 = new("./seq_loop_status20.csv");
    seq_loop_monitor_20 = new(seq_loop_intf_20,seq_loop_csv_dumper_20);
    seq_loop_csv_dumper_21 = new("./seq_loop_status21.csv");
    seq_loop_monitor_21 = new(seq_loop_intf_21,seq_loop_csv_dumper_21);
    seq_loop_csv_dumper_22 = new("./seq_loop_status22.csv");
    seq_loop_monitor_22 = new(seq_loop_intf_22,seq_loop_csv_dumper_22);
    seq_loop_csv_dumper_23 = new("./seq_loop_status23.csv");
    seq_loop_monitor_23 = new(seq_loop_intf_23,seq_loop_csv_dumper_23);
    seq_loop_csv_dumper_24 = new("./seq_loop_status24.csv");
    seq_loop_monitor_24 = new(seq_loop_intf_24,seq_loop_csv_dumper_24);
    seq_loop_csv_dumper_25 = new("./seq_loop_status25.csv");
    seq_loop_monitor_25 = new(seq_loop_intf_25,seq_loop_csv_dumper_25);
    seq_loop_csv_dumper_26 = new("./seq_loop_status26.csv");
    seq_loop_monitor_26 = new(seq_loop_intf_26,seq_loop_csv_dumper_26);
    seq_loop_csv_dumper_27 = new("./seq_loop_status27.csv");
    seq_loop_monitor_27 = new(seq_loop_intf_27,seq_loop_csv_dumper_27);
    seq_loop_csv_dumper_28 = new("./seq_loop_status28.csv");
    seq_loop_monitor_28 = new(seq_loop_intf_28,seq_loop_csv_dumper_28);
    seq_loop_csv_dumper_29 = new("./seq_loop_status29.csv");
    seq_loop_monitor_29 = new(seq_loop_intf_29,seq_loop_csv_dumper_29);
    seq_loop_csv_dumper_30 = new("./seq_loop_status30.csv");
    seq_loop_monitor_30 = new(seq_loop_intf_30,seq_loop_csv_dumper_30);
    seq_loop_csv_dumper_31 = new("./seq_loop_status31.csv");
    seq_loop_monitor_31 = new(seq_loop_intf_31,seq_loop_csv_dumper_31);
    seq_loop_csv_dumper_32 = new("./seq_loop_status32.csv");
    seq_loop_monitor_32 = new(seq_loop_intf_32,seq_loop_csv_dumper_32);
    seq_loop_csv_dumper_33 = new("./seq_loop_status33.csv");
    seq_loop_monitor_33 = new(seq_loop_intf_33,seq_loop_csv_dumper_33);
    seq_loop_csv_dumper_34 = new("./seq_loop_status34.csv");
    seq_loop_monitor_34 = new(seq_loop_intf_34,seq_loop_csv_dumper_34);
    seq_loop_csv_dumper_35 = new("./seq_loop_status35.csv");
    seq_loop_monitor_35 = new(seq_loop_intf_35,seq_loop_csv_dumper_35);
    seq_loop_csv_dumper_36 = new("./seq_loop_status36.csv");
    seq_loop_monitor_36 = new(seq_loop_intf_36,seq_loop_csv_dumper_36);
    seq_loop_csv_dumper_37 = new("./seq_loop_status37.csv");
    seq_loop_monitor_37 = new(seq_loop_intf_37,seq_loop_csv_dumper_37);
    seq_loop_csv_dumper_38 = new("./seq_loop_status38.csv");
    seq_loop_monitor_38 = new(seq_loop_intf_38,seq_loop_csv_dumper_38);
    seq_loop_csv_dumper_39 = new("./seq_loop_status39.csv");
    seq_loop_monitor_39 = new(seq_loop_intf_39,seq_loop_csv_dumper_39);
    seq_loop_csv_dumper_40 = new("./seq_loop_status40.csv");
    seq_loop_monitor_40 = new(seq_loop_intf_40,seq_loop_csv_dumper_40);
    seq_loop_csv_dumper_41 = new("./seq_loop_status41.csv");
    seq_loop_monitor_41 = new(seq_loop_intf_41,seq_loop_csv_dumper_41);
    seq_loop_csv_dumper_42 = new("./seq_loop_status42.csv");
    seq_loop_monitor_42 = new(seq_loop_intf_42,seq_loop_csv_dumper_42);
    seq_loop_csv_dumper_43 = new("./seq_loop_status43.csv");
    seq_loop_monitor_43 = new(seq_loop_intf_43,seq_loop_csv_dumper_43);
    seq_loop_csv_dumper_44 = new("./seq_loop_status44.csv");
    seq_loop_monitor_44 = new(seq_loop_intf_44,seq_loop_csv_dumper_44);
    seq_loop_csv_dumper_45 = new("./seq_loop_status45.csv");
    seq_loop_monitor_45 = new(seq_loop_intf_45,seq_loop_csv_dumper_45);
    seq_loop_csv_dumper_46 = new("./seq_loop_status46.csv");
    seq_loop_monitor_46 = new(seq_loop_intf_46,seq_loop_csv_dumper_46);
    seq_loop_csv_dumper_47 = new("./seq_loop_status47.csv");
    seq_loop_monitor_47 = new(seq_loop_intf_47,seq_loop_csv_dumper_47);
    seq_loop_csv_dumper_48 = new("./seq_loop_status48.csv");
    seq_loop_monitor_48 = new(seq_loop_intf_48,seq_loop_csv_dumper_48);
    seq_loop_csv_dumper_49 = new("./seq_loop_status49.csv");
    seq_loop_monitor_49 = new(seq_loop_intf_49,seq_loop_csv_dumper_49);
    seq_loop_csv_dumper_50 = new("./seq_loop_status50.csv");
    seq_loop_monitor_50 = new(seq_loop_intf_50,seq_loop_csv_dumper_50);
    seq_loop_csv_dumper_51 = new("./seq_loop_status51.csv");
    seq_loop_monitor_51 = new(seq_loop_intf_51,seq_loop_csv_dumper_51);
    seq_loop_csv_dumper_52 = new("./seq_loop_status52.csv");
    seq_loop_monitor_52 = new(seq_loop_intf_52,seq_loop_csv_dumper_52);
    seq_loop_csv_dumper_53 = new("./seq_loop_status53.csv");
    seq_loop_monitor_53 = new(seq_loop_intf_53,seq_loop_csv_dumper_53);
    seq_loop_csv_dumper_54 = new("./seq_loop_status54.csv");
    seq_loop_monitor_54 = new(seq_loop_intf_54,seq_loop_csv_dumper_54);
    seq_loop_csv_dumper_55 = new("./seq_loop_status55.csv");
    seq_loop_monitor_55 = new(seq_loop_intf_55,seq_loop_csv_dumper_55);
    seq_loop_csv_dumper_56 = new("./seq_loop_status56.csv");
    seq_loop_monitor_56 = new(seq_loop_intf_56,seq_loop_csv_dumper_56);
    seq_loop_csv_dumper_57 = new("./seq_loop_status57.csv");
    seq_loop_monitor_57 = new(seq_loop_intf_57,seq_loop_csv_dumper_57);
    seq_loop_csv_dumper_58 = new("./seq_loop_status58.csv");
    seq_loop_monitor_58 = new(seq_loop_intf_58,seq_loop_csv_dumper_58);
    seq_loop_csv_dumper_59 = new("./seq_loop_status59.csv");
    seq_loop_monitor_59 = new(seq_loop_intf_59,seq_loop_csv_dumper_59);
    seq_loop_csv_dumper_60 = new("./seq_loop_status60.csv");
    seq_loop_monitor_60 = new(seq_loop_intf_60,seq_loop_csv_dumper_60);
    seq_loop_csv_dumper_61 = new("./seq_loop_status61.csv");
    seq_loop_monitor_61 = new(seq_loop_intf_61,seq_loop_csv_dumper_61);
    seq_loop_csv_dumper_62 = new("./seq_loop_status62.csv");
    seq_loop_monitor_62 = new(seq_loop_intf_62,seq_loop_csv_dumper_62);
    seq_loop_csv_dumper_63 = new("./seq_loop_status63.csv");
    seq_loop_monitor_63 = new(seq_loop_intf_63,seq_loop_csv_dumper_63);
    seq_loop_csv_dumper_64 = new("./seq_loop_status64.csv");
    seq_loop_monitor_64 = new(seq_loop_intf_64,seq_loop_csv_dumper_64);
    seq_loop_csv_dumper_65 = new("./seq_loop_status65.csv");
    seq_loop_monitor_65 = new(seq_loop_intf_65,seq_loop_csv_dumper_65);
    seq_loop_csv_dumper_66 = new("./seq_loop_status66.csv");
    seq_loop_monitor_66 = new(seq_loop_intf_66,seq_loop_csv_dumper_66);
    seq_loop_csv_dumper_67 = new("./seq_loop_status67.csv");
    seq_loop_monitor_67 = new(seq_loop_intf_67,seq_loop_csv_dumper_67);
    seq_loop_csv_dumper_68 = new("./seq_loop_status68.csv");
    seq_loop_monitor_68 = new(seq_loop_intf_68,seq_loop_csv_dumper_68);
    seq_loop_csv_dumper_69 = new("./seq_loop_status69.csv");
    seq_loop_monitor_69 = new(seq_loop_intf_69,seq_loop_csv_dumper_69);
    seq_loop_csv_dumper_70 = new("./seq_loop_status70.csv");
    seq_loop_monitor_70 = new(seq_loop_intf_70,seq_loop_csv_dumper_70);
    seq_loop_csv_dumper_71 = new("./seq_loop_status71.csv");
    seq_loop_monitor_71 = new(seq_loop_intf_71,seq_loop_csv_dumper_71);
    seq_loop_csv_dumper_72 = new("./seq_loop_status72.csv");
    seq_loop_monitor_72 = new(seq_loop_intf_72,seq_loop_csv_dumper_72);
    seq_loop_csv_dumper_73 = new("./seq_loop_status73.csv");
    seq_loop_monitor_73 = new(seq_loop_intf_73,seq_loop_csv_dumper_73);
    seq_loop_csv_dumper_74 = new("./seq_loop_status74.csv");
    seq_loop_monitor_74 = new(seq_loop_intf_74,seq_loop_csv_dumper_74);
    seq_loop_csv_dumper_75 = new("./seq_loop_status75.csv");
    seq_loop_monitor_75 = new(seq_loop_intf_75,seq_loop_csv_dumper_75);
    seq_loop_csv_dumper_76 = new("./seq_loop_status76.csv");
    seq_loop_monitor_76 = new(seq_loop_intf_76,seq_loop_csv_dumper_76);
    seq_loop_csv_dumper_77 = new("./seq_loop_status77.csv");
    seq_loop_monitor_77 = new(seq_loop_intf_77,seq_loop_csv_dumper_77);
    seq_loop_csv_dumper_78 = new("./seq_loop_status78.csv");
    seq_loop_monitor_78 = new(seq_loop_intf_78,seq_loop_csv_dumper_78);
    seq_loop_csv_dumper_79 = new("./seq_loop_status79.csv");
    seq_loop_monitor_79 = new(seq_loop_intf_79,seq_loop_csv_dumper_79);
    seq_loop_csv_dumper_80 = new("./seq_loop_status80.csv");
    seq_loop_monitor_80 = new(seq_loop_intf_80,seq_loop_csv_dumper_80);
    seq_loop_csv_dumper_81 = new("./seq_loop_status81.csv");
    seq_loop_monitor_81 = new(seq_loop_intf_81,seq_loop_csv_dumper_81);
    seq_loop_csv_dumper_82 = new("./seq_loop_status82.csv");
    seq_loop_monitor_82 = new(seq_loop_intf_82,seq_loop_csv_dumper_82);
    seq_loop_csv_dumper_83 = new("./seq_loop_status83.csv");
    seq_loop_monitor_83 = new(seq_loop_intf_83,seq_loop_csv_dumper_83);
    seq_loop_csv_dumper_84 = new("./seq_loop_status84.csv");
    seq_loop_monitor_84 = new(seq_loop_intf_84,seq_loop_csv_dumper_84);
    seq_loop_csv_dumper_85 = new("./seq_loop_status85.csv");
    seq_loop_monitor_85 = new(seq_loop_intf_85,seq_loop_csv_dumper_85);
    seq_loop_csv_dumper_86 = new("./seq_loop_status86.csv");
    seq_loop_monitor_86 = new(seq_loop_intf_86,seq_loop_csv_dumper_86);
    seq_loop_csv_dumper_87 = new("./seq_loop_status87.csv");
    seq_loop_monitor_87 = new(seq_loop_intf_87,seq_loop_csv_dumper_87);
    seq_loop_csv_dumper_88 = new("./seq_loop_status88.csv");
    seq_loop_monitor_88 = new(seq_loop_intf_88,seq_loop_csv_dumper_88);
    seq_loop_csv_dumper_89 = new("./seq_loop_status89.csv");
    seq_loop_monitor_89 = new(seq_loop_intf_89,seq_loop_csv_dumper_89);
    seq_loop_csv_dumper_90 = new("./seq_loop_status90.csv");
    seq_loop_monitor_90 = new(seq_loop_intf_90,seq_loop_csv_dumper_90);
    seq_loop_csv_dumper_91 = new("./seq_loop_status91.csv");
    seq_loop_monitor_91 = new(seq_loop_intf_91,seq_loop_csv_dumper_91);
    seq_loop_csv_dumper_92 = new("./seq_loop_status92.csv");
    seq_loop_monitor_92 = new(seq_loop_intf_92,seq_loop_csv_dumper_92);
    seq_loop_csv_dumper_93 = new("./seq_loop_status93.csv");
    seq_loop_monitor_93 = new(seq_loop_intf_93,seq_loop_csv_dumper_93);
    seq_loop_csv_dumper_94 = new("./seq_loop_status94.csv");
    seq_loop_monitor_94 = new(seq_loop_intf_94,seq_loop_csv_dumper_94);
    seq_loop_csv_dumper_95 = new("./seq_loop_status95.csv");
    seq_loop_monitor_95 = new(seq_loop_intf_95,seq_loop_csv_dumper_95);
    seq_loop_csv_dumper_96 = new("./seq_loop_status96.csv");
    seq_loop_monitor_96 = new(seq_loop_intf_96,seq_loop_csv_dumper_96);
    seq_loop_csv_dumper_97 = new("./seq_loop_status97.csv");
    seq_loop_monitor_97 = new(seq_loop_intf_97,seq_loop_csv_dumper_97);
    seq_loop_csv_dumper_98 = new("./seq_loop_status98.csv");
    seq_loop_monitor_98 = new(seq_loop_intf_98,seq_loop_csv_dumper_98);
    seq_loop_csv_dumper_99 = new("./seq_loop_status99.csv");
    seq_loop_monitor_99 = new(seq_loop_intf_99,seq_loop_csv_dumper_99);
    seq_loop_csv_dumper_100 = new("./seq_loop_status100.csv");
    seq_loop_monitor_100 = new(seq_loop_intf_100,seq_loop_csv_dumper_100);
    seq_loop_csv_dumper_101 = new("./seq_loop_status101.csv");
    seq_loop_monitor_101 = new(seq_loop_intf_101,seq_loop_csv_dumper_101);
    seq_loop_csv_dumper_102 = new("./seq_loop_status102.csv");
    seq_loop_monitor_102 = new(seq_loop_intf_102,seq_loop_csv_dumper_102);
    seq_loop_csv_dumper_103 = new("./seq_loop_status103.csv");
    seq_loop_monitor_103 = new(seq_loop_intf_103,seq_loop_csv_dumper_103);
    seq_loop_csv_dumper_104 = new("./seq_loop_status104.csv");
    seq_loop_monitor_104 = new(seq_loop_intf_104,seq_loop_csv_dumper_104);
    seq_loop_csv_dumper_105 = new("./seq_loop_status105.csv");
    seq_loop_monitor_105 = new(seq_loop_intf_105,seq_loop_csv_dumper_105);
    seq_loop_csv_dumper_106 = new("./seq_loop_status106.csv");
    seq_loop_monitor_106 = new(seq_loop_intf_106,seq_loop_csv_dumper_106);
    seq_loop_csv_dumper_107 = new("./seq_loop_status107.csv");
    seq_loop_monitor_107 = new(seq_loop_intf_107,seq_loop_csv_dumper_107);
    seq_loop_csv_dumper_108 = new("./seq_loop_status108.csv");
    seq_loop_monitor_108 = new(seq_loop_intf_108,seq_loop_csv_dumper_108);
    seq_loop_csv_dumper_109 = new("./seq_loop_status109.csv");
    seq_loop_monitor_109 = new(seq_loop_intf_109,seq_loop_csv_dumper_109);
    seq_loop_csv_dumper_110 = new("./seq_loop_status110.csv");
    seq_loop_monitor_110 = new(seq_loop_intf_110,seq_loop_csv_dumper_110);
    seq_loop_csv_dumper_111 = new("./seq_loop_status111.csv");
    seq_loop_monitor_111 = new(seq_loop_intf_111,seq_loop_csv_dumper_111);
    seq_loop_csv_dumper_112 = new("./seq_loop_status112.csv");
    seq_loop_monitor_112 = new(seq_loop_intf_112,seq_loop_csv_dumper_112);
    seq_loop_csv_dumper_113 = new("./seq_loop_status113.csv");
    seq_loop_monitor_113 = new(seq_loop_intf_113,seq_loop_csv_dumper_113);
    seq_loop_csv_dumper_114 = new("./seq_loop_status114.csv");
    seq_loop_monitor_114 = new(seq_loop_intf_114,seq_loop_csv_dumper_114);
    seq_loop_csv_dumper_115 = new("./seq_loop_status115.csv");
    seq_loop_monitor_115 = new(seq_loop_intf_115,seq_loop_csv_dumper_115);
    seq_loop_csv_dumper_116 = new("./seq_loop_status116.csv");
    seq_loop_monitor_116 = new(seq_loop_intf_116,seq_loop_csv_dumper_116);
    seq_loop_csv_dumper_117 = new("./seq_loop_status117.csv");
    seq_loop_monitor_117 = new(seq_loop_intf_117,seq_loop_csv_dumper_117);
    seq_loop_csv_dumper_118 = new("./seq_loop_status118.csv");
    seq_loop_monitor_118 = new(seq_loop_intf_118,seq_loop_csv_dumper_118);
    seq_loop_csv_dumper_119 = new("./seq_loop_status119.csv");
    seq_loop_monitor_119 = new(seq_loop_intf_119,seq_loop_csv_dumper_119);
    seq_loop_csv_dumper_120 = new("./seq_loop_status120.csv");
    seq_loop_monitor_120 = new(seq_loop_intf_120,seq_loop_csv_dumper_120);
    seq_loop_csv_dumper_121 = new("./seq_loop_status121.csv");
    seq_loop_monitor_121 = new(seq_loop_intf_121,seq_loop_csv_dumper_121);
    seq_loop_csv_dumper_122 = new("./seq_loop_status122.csv");
    seq_loop_monitor_122 = new(seq_loop_intf_122,seq_loop_csv_dumper_122);
    seq_loop_csv_dumper_123 = new("./seq_loop_status123.csv");
    seq_loop_monitor_123 = new(seq_loop_intf_123,seq_loop_csv_dumper_123);
    seq_loop_csv_dumper_124 = new("./seq_loop_status124.csv");
    seq_loop_monitor_124 = new(seq_loop_intf_124,seq_loop_csv_dumper_124);
    seq_loop_csv_dumper_125 = new("./seq_loop_status125.csv");
    seq_loop_monitor_125 = new(seq_loop_intf_125,seq_loop_csv_dumper_125);
    seq_loop_csv_dumper_126 = new("./seq_loop_status126.csv");
    seq_loop_monitor_126 = new(seq_loop_intf_126,seq_loop_csv_dumper_126);
    seq_loop_csv_dumper_127 = new("./seq_loop_status127.csv");
    seq_loop_monitor_127 = new(seq_loop_intf_127,seq_loop_csv_dumper_127);
    seq_loop_csv_dumper_128 = new("./seq_loop_status128.csv");
    seq_loop_monitor_128 = new(seq_loop_intf_128,seq_loop_csv_dumper_128);
    seq_loop_csv_dumper_129 = new("./seq_loop_status129.csv");
    seq_loop_monitor_129 = new(seq_loop_intf_129,seq_loop_csv_dumper_129);
    seq_loop_csv_dumper_130 = new("./seq_loop_status130.csv");
    seq_loop_monitor_130 = new(seq_loop_intf_130,seq_loop_csv_dumper_130);
    seq_loop_csv_dumper_131 = new("./seq_loop_status131.csv");
    seq_loop_monitor_131 = new(seq_loop_intf_131,seq_loop_csv_dumper_131);
    seq_loop_csv_dumper_132 = new("./seq_loop_status132.csv");
    seq_loop_monitor_132 = new(seq_loop_intf_132,seq_loop_csv_dumper_132);
    seq_loop_csv_dumper_133 = new("./seq_loop_status133.csv");
    seq_loop_monitor_133 = new(seq_loop_intf_133,seq_loop_csv_dumper_133);
    seq_loop_csv_dumper_134 = new("./seq_loop_status134.csv");
    seq_loop_monitor_134 = new(seq_loop_intf_134,seq_loop_csv_dumper_134);
    seq_loop_csv_dumper_135 = new("./seq_loop_status135.csv");
    seq_loop_monitor_135 = new(seq_loop_intf_135,seq_loop_csv_dumper_135);
    seq_loop_csv_dumper_136 = new("./seq_loop_status136.csv");
    seq_loop_monitor_136 = new(seq_loop_intf_136,seq_loop_csv_dumper_136);
    seq_loop_csv_dumper_137 = new("./seq_loop_status137.csv");
    seq_loop_monitor_137 = new(seq_loop_intf_137,seq_loop_csv_dumper_137);
    seq_loop_csv_dumper_138 = new("./seq_loop_status138.csv");
    seq_loop_monitor_138 = new(seq_loop_intf_138,seq_loop_csv_dumper_138);
    seq_loop_csv_dumper_139 = new("./seq_loop_status139.csv");
    seq_loop_monitor_139 = new(seq_loop_intf_139,seq_loop_csv_dumper_139);
    seq_loop_csv_dumper_140 = new("./seq_loop_status140.csv");
    seq_loop_monitor_140 = new(seq_loop_intf_140,seq_loop_csv_dumper_140);
    seq_loop_csv_dumper_141 = new("./seq_loop_status141.csv");
    seq_loop_monitor_141 = new(seq_loop_intf_141,seq_loop_csv_dumper_141);
    seq_loop_csv_dumper_142 = new("./seq_loop_status142.csv");
    seq_loop_monitor_142 = new(seq_loop_intf_142,seq_loop_csv_dumper_142);
    seq_loop_csv_dumper_143 = new("./seq_loop_status143.csv");
    seq_loop_monitor_143 = new(seq_loop_intf_143,seq_loop_csv_dumper_143);
    seq_loop_csv_dumper_144 = new("./seq_loop_status144.csv");
    seq_loop_monitor_144 = new(seq_loop_intf_144,seq_loop_csv_dumper_144);
    seq_loop_csv_dumper_145 = new("./seq_loop_status145.csv");
    seq_loop_monitor_145 = new(seq_loop_intf_145,seq_loop_csv_dumper_145);
    seq_loop_csv_dumper_146 = new("./seq_loop_status146.csv");
    seq_loop_monitor_146 = new(seq_loop_intf_146,seq_loop_csv_dumper_146);
    seq_loop_csv_dumper_147 = new("./seq_loop_status147.csv");
    seq_loop_monitor_147 = new(seq_loop_intf_147,seq_loop_csv_dumper_147);
    seq_loop_csv_dumper_148 = new("./seq_loop_status148.csv");
    seq_loop_monitor_148 = new(seq_loop_intf_148,seq_loop_csv_dumper_148);
    seq_loop_csv_dumper_149 = new("./seq_loop_status149.csv");
    seq_loop_monitor_149 = new(seq_loop_intf_149,seq_loop_csv_dumper_149);
    seq_loop_csv_dumper_150 = new("./seq_loop_status150.csv");
    seq_loop_monitor_150 = new(seq_loop_intf_150,seq_loop_csv_dumper_150);
    seq_loop_csv_dumper_151 = new("./seq_loop_status151.csv");
    seq_loop_monitor_151 = new(seq_loop_intf_151,seq_loop_csv_dumper_151);
    seq_loop_csv_dumper_152 = new("./seq_loop_status152.csv");
    seq_loop_monitor_152 = new(seq_loop_intf_152,seq_loop_csv_dumper_152);
    seq_loop_csv_dumper_153 = new("./seq_loop_status153.csv");
    seq_loop_monitor_153 = new(seq_loop_intf_153,seq_loop_csv_dumper_153);
    seq_loop_csv_dumper_154 = new("./seq_loop_status154.csv");
    seq_loop_monitor_154 = new(seq_loop_intf_154,seq_loop_csv_dumper_154);
    seq_loop_csv_dumper_155 = new("./seq_loop_status155.csv");
    seq_loop_monitor_155 = new(seq_loop_intf_155,seq_loop_csv_dumper_155);
    seq_loop_csv_dumper_156 = new("./seq_loop_status156.csv");
    seq_loop_monitor_156 = new(seq_loop_intf_156,seq_loop_csv_dumper_156);
    seq_loop_csv_dumper_157 = new("./seq_loop_status157.csv");
    seq_loop_monitor_157 = new(seq_loop_intf_157,seq_loop_csv_dumper_157);
    seq_loop_csv_dumper_158 = new("./seq_loop_status158.csv");
    seq_loop_monitor_158 = new(seq_loop_intf_158,seq_loop_csv_dumper_158);
    seq_loop_csv_dumper_159 = new("./seq_loop_status159.csv");
    seq_loop_monitor_159 = new(seq_loop_intf_159,seq_loop_csv_dumper_159);
    seq_loop_csv_dumper_160 = new("./seq_loop_status160.csv");
    seq_loop_monitor_160 = new(seq_loop_intf_160,seq_loop_csv_dumper_160);
    seq_loop_csv_dumper_161 = new("./seq_loop_status161.csv");
    seq_loop_monitor_161 = new(seq_loop_intf_161,seq_loop_csv_dumper_161);
    seq_loop_csv_dumper_162 = new("./seq_loop_status162.csv");
    seq_loop_monitor_162 = new(seq_loop_intf_162,seq_loop_csv_dumper_162);
    seq_loop_csv_dumper_163 = new("./seq_loop_status163.csv");
    seq_loop_monitor_163 = new(seq_loop_intf_163,seq_loop_csv_dumper_163);
    seq_loop_csv_dumper_164 = new("./seq_loop_status164.csv");
    seq_loop_monitor_164 = new(seq_loop_intf_164,seq_loop_csv_dumper_164);
    seq_loop_csv_dumper_165 = new("./seq_loop_status165.csv");
    seq_loop_monitor_165 = new(seq_loop_intf_165,seq_loop_csv_dumper_165);
    seq_loop_csv_dumper_166 = new("./seq_loop_status166.csv");
    seq_loop_monitor_166 = new(seq_loop_intf_166,seq_loop_csv_dumper_166);
    seq_loop_csv_dumper_167 = new("./seq_loop_status167.csv");
    seq_loop_monitor_167 = new(seq_loop_intf_167,seq_loop_csv_dumper_167);
    seq_loop_csv_dumper_168 = new("./seq_loop_status168.csv");
    seq_loop_monitor_168 = new(seq_loop_intf_168,seq_loop_csv_dumper_168);
    seq_loop_csv_dumper_169 = new("./seq_loop_status169.csv");
    seq_loop_monitor_169 = new(seq_loop_intf_169,seq_loop_csv_dumper_169);
    seq_loop_csv_dumper_170 = new("./seq_loop_status170.csv");
    seq_loop_monitor_170 = new(seq_loop_intf_170,seq_loop_csv_dumper_170);
    seq_loop_csv_dumper_171 = new("./seq_loop_status171.csv");
    seq_loop_monitor_171 = new(seq_loop_intf_171,seq_loop_csv_dumper_171);
    seq_loop_csv_dumper_172 = new("./seq_loop_status172.csv");
    seq_loop_monitor_172 = new(seq_loop_intf_172,seq_loop_csv_dumper_172);
    seq_loop_csv_dumper_173 = new("./seq_loop_status173.csv");
    seq_loop_monitor_173 = new(seq_loop_intf_173,seq_loop_csv_dumper_173);
    seq_loop_csv_dumper_174 = new("./seq_loop_status174.csv");
    seq_loop_monitor_174 = new(seq_loop_intf_174,seq_loop_csv_dumper_174);
    seq_loop_csv_dumper_175 = new("./seq_loop_status175.csv");
    seq_loop_monitor_175 = new(seq_loop_intf_175,seq_loop_csv_dumper_175);
    seq_loop_csv_dumper_176 = new("./seq_loop_status176.csv");
    seq_loop_monitor_176 = new(seq_loop_intf_176,seq_loop_csv_dumper_176);
    seq_loop_csv_dumper_177 = new("./seq_loop_status177.csv");
    seq_loop_monitor_177 = new(seq_loop_intf_177,seq_loop_csv_dumper_177);
    seq_loop_csv_dumper_178 = new("./seq_loop_status178.csv");
    seq_loop_monitor_178 = new(seq_loop_intf_178,seq_loop_csv_dumper_178);
    seq_loop_csv_dumper_179 = new("./seq_loop_status179.csv");
    seq_loop_monitor_179 = new(seq_loop_intf_179,seq_loop_csv_dumper_179);
    seq_loop_csv_dumper_180 = new("./seq_loop_status180.csv");
    seq_loop_monitor_180 = new(seq_loop_intf_180,seq_loop_csv_dumper_180);
    seq_loop_csv_dumper_181 = new("./seq_loop_status181.csv");
    seq_loop_monitor_181 = new(seq_loop_intf_181,seq_loop_csv_dumper_181);
    seq_loop_csv_dumper_182 = new("./seq_loop_status182.csv");
    seq_loop_monitor_182 = new(seq_loop_intf_182,seq_loop_csv_dumper_182);
    seq_loop_csv_dumper_183 = new("./seq_loop_status183.csv");
    seq_loop_monitor_183 = new(seq_loop_intf_183,seq_loop_csv_dumper_183);
    seq_loop_csv_dumper_184 = new("./seq_loop_status184.csv");
    seq_loop_monitor_184 = new(seq_loop_intf_184,seq_loop_csv_dumper_184);
    seq_loop_csv_dumper_185 = new("./seq_loop_status185.csv");
    seq_loop_monitor_185 = new(seq_loop_intf_185,seq_loop_csv_dumper_185);
    seq_loop_csv_dumper_186 = new("./seq_loop_status186.csv");
    seq_loop_monitor_186 = new(seq_loop_intf_186,seq_loop_csv_dumper_186);
    seq_loop_csv_dumper_187 = new("./seq_loop_status187.csv");
    seq_loop_monitor_187 = new(seq_loop_intf_187,seq_loop_csv_dumper_187);
    seq_loop_csv_dumper_188 = new("./seq_loop_status188.csv");
    seq_loop_monitor_188 = new(seq_loop_intf_188,seq_loop_csv_dumper_188);
    seq_loop_csv_dumper_189 = new("./seq_loop_status189.csv");
    seq_loop_monitor_189 = new(seq_loop_intf_189,seq_loop_csv_dumper_189);
    seq_loop_csv_dumper_190 = new("./seq_loop_status190.csv");
    seq_loop_monitor_190 = new(seq_loop_intf_190,seq_loop_csv_dumper_190);
    seq_loop_csv_dumper_191 = new("./seq_loop_status191.csv");
    seq_loop_monitor_191 = new(seq_loop_intf_191,seq_loop_csv_dumper_191);
    seq_loop_csv_dumper_192 = new("./seq_loop_status192.csv");
    seq_loop_monitor_192 = new(seq_loop_intf_192,seq_loop_csv_dumper_192);
    seq_loop_csv_dumper_193 = new("./seq_loop_status193.csv");
    seq_loop_monitor_193 = new(seq_loop_intf_193,seq_loop_csv_dumper_193);
    seq_loop_csv_dumper_194 = new("./seq_loop_status194.csv");
    seq_loop_monitor_194 = new(seq_loop_intf_194,seq_loop_csv_dumper_194);
    seq_loop_csv_dumper_195 = new("./seq_loop_status195.csv");
    seq_loop_monitor_195 = new(seq_loop_intf_195,seq_loop_csv_dumper_195);
    seq_loop_csv_dumper_196 = new("./seq_loop_status196.csv");
    seq_loop_monitor_196 = new(seq_loop_intf_196,seq_loop_csv_dumper_196);
    seq_loop_csv_dumper_197 = new("./seq_loop_status197.csv");
    seq_loop_monitor_197 = new(seq_loop_intf_197,seq_loop_csv_dumper_197);
    seq_loop_csv_dumper_198 = new("./seq_loop_status198.csv");
    seq_loop_monitor_198 = new(seq_loop_intf_198,seq_loop_csv_dumper_198);
    seq_loop_csv_dumper_199 = new("./seq_loop_status199.csv");
    seq_loop_monitor_199 = new(seq_loop_intf_199,seq_loop_csv_dumper_199);
    seq_loop_csv_dumper_200 = new("./seq_loop_status200.csv");
    seq_loop_monitor_200 = new(seq_loop_intf_200,seq_loop_csv_dumper_200);
    seq_loop_csv_dumper_201 = new("./seq_loop_status201.csv");
    seq_loop_monitor_201 = new(seq_loop_intf_201,seq_loop_csv_dumper_201);
    seq_loop_csv_dumper_202 = new("./seq_loop_status202.csv");
    seq_loop_monitor_202 = new(seq_loop_intf_202,seq_loop_csv_dumper_202);
    seq_loop_csv_dumper_203 = new("./seq_loop_status203.csv");
    seq_loop_monitor_203 = new(seq_loop_intf_203,seq_loop_csv_dumper_203);
    seq_loop_csv_dumper_204 = new("./seq_loop_status204.csv");
    seq_loop_monitor_204 = new(seq_loop_intf_204,seq_loop_csv_dumper_204);
    seq_loop_csv_dumper_205 = new("./seq_loop_status205.csv");
    seq_loop_monitor_205 = new(seq_loop_intf_205,seq_loop_csv_dumper_205);
    seq_loop_csv_dumper_206 = new("./seq_loop_status206.csv");
    seq_loop_monitor_206 = new(seq_loop_intf_206,seq_loop_csv_dumper_206);
    seq_loop_csv_dumper_207 = new("./seq_loop_status207.csv");
    seq_loop_monitor_207 = new(seq_loop_intf_207,seq_loop_csv_dumper_207);
    seq_loop_csv_dumper_208 = new("./seq_loop_status208.csv");
    seq_loop_monitor_208 = new(seq_loop_intf_208,seq_loop_csv_dumper_208);
    seq_loop_csv_dumper_209 = new("./seq_loop_status209.csv");
    seq_loop_monitor_209 = new(seq_loop_intf_209,seq_loop_csv_dumper_209);
    seq_loop_csv_dumper_210 = new("./seq_loop_status210.csv");
    seq_loop_monitor_210 = new(seq_loop_intf_210,seq_loop_csv_dumper_210);
    seq_loop_csv_dumper_211 = new("./seq_loop_status211.csv");
    seq_loop_monitor_211 = new(seq_loop_intf_211,seq_loop_csv_dumper_211);
    seq_loop_csv_dumper_212 = new("./seq_loop_status212.csv");
    seq_loop_monitor_212 = new(seq_loop_intf_212,seq_loop_csv_dumper_212);
    seq_loop_csv_dumper_213 = new("./seq_loop_status213.csv");
    seq_loop_monitor_213 = new(seq_loop_intf_213,seq_loop_csv_dumper_213);
    seq_loop_csv_dumper_214 = new("./seq_loop_status214.csv");
    seq_loop_monitor_214 = new(seq_loop_intf_214,seq_loop_csv_dumper_214);
    seq_loop_csv_dumper_215 = new("./seq_loop_status215.csv");
    seq_loop_monitor_215 = new(seq_loop_intf_215,seq_loop_csv_dumper_215);
    seq_loop_csv_dumper_216 = new("./seq_loop_status216.csv");
    seq_loop_monitor_216 = new(seq_loop_intf_216,seq_loop_csv_dumper_216);
    seq_loop_csv_dumper_217 = new("./seq_loop_status217.csv");
    seq_loop_monitor_217 = new(seq_loop_intf_217,seq_loop_csv_dumper_217);
    seq_loop_csv_dumper_218 = new("./seq_loop_status218.csv");
    seq_loop_monitor_218 = new(seq_loop_intf_218,seq_loop_csv_dumper_218);
    seq_loop_csv_dumper_219 = new("./seq_loop_status219.csv");
    seq_loop_monitor_219 = new(seq_loop_intf_219,seq_loop_csv_dumper_219);
    seq_loop_csv_dumper_220 = new("./seq_loop_status220.csv");
    seq_loop_monitor_220 = new(seq_loop_intf_220,seq_loop_csv_dumper_220);
    seq_loop_csv_dumper_221 = new("./seq_loop_status221.csv");
    seq_loop_monitor_221 = new(seq_loop_intf_221,seq_loop_csv_dumper_221);
    seq_loop_csv_dumper_222 = new("./seq_loop_status222.csv");
    seq_loop_monitor_222 = new(seq_loop_intf_222,seq_loop_csv_dumper_222);
    seq_loop_csv_dumper_223 = new("./seq_loop_status223.csv");
    seq_loop_monitor_223 = new(seq_loop_intf_223,seq_loop_csv_dumper_223);
    seq_loop_csv_dumper_224 = new("./seq_loop_status224.csv");
    seq_loop_monitor_224 = new(seq_loop_intf_224,seq_loop_csv_dumper_224);
    seq_loop_csv_dumper_225 = new("./seq_loop_status225.csv");
    seq_loop_monitor_225 = new(seq_loop_intf_225,seq_loop_csv_dumper_225);
    seq_loop_csv_dumper_226 = new("./seq_loop_status226.csv");
    seq_loop_monitor_226 = new(seq_loop_intf_226,seq_loop_csv_dumper_226);
    seq_loop_csv_dumper_227 = new("./seq_loop_status227.csv");
    seq_loop_monitor_227 = new(seq_loop_intf_227,seq_loop_csv_dumper_227);
    seq_loop_csv_dumper_228 = new("./seq_loop_status228.csv");
    seq_loop_monitor_228 = new(seq_loop_intf_228,seq_loop_csv_dumper_228);
    seq_loop_csv_dumper_229 = new("./seq_loop_status229.csv");
    seq_loop_monitor_229 = new(seq_loop_intf_229,seq_loop_csv_dumper_229);
    seq_loop_csv_dumper_230 = new("./seq_loop_status230.csv");
    seq_loop_monitor_230 = new(seq_loop_intf_230,seq_loop_csv_dumper_230);
    seq_loop_csv_dumper_231 = new("./seq_loop_status231.csv");
    seq_loop_monitor_231 = new(seq_loop_intf_231,seq_loop_csv_dumper_231);
    seq_loop_csv_dumper_232 = new("./seq_loop_status232.csv");
    seq_loop_monitor_232 = new(seq_loop_intf_232,seq_loop_csv_dumper_232);
    seq_loop_csv_dumper_233 = new("./seq_loop_status233.csv");
    seq_loop_monitor_233 = new(seq_loop_intf_233,seq_loop_csv_dumper_233);
    seq_loop_csv_dumper_234 = new("./seq_loop_status234.csv");
    seq_loop_monitor_234 = new(seq_loop_intf_234,seq_loop_csv_dumper_234);
    seq_loop_csv_dumper_235 = new("./seq_loop_status235.csv");
    seq_loop_monitor_235 = new(seq_loop_intf_235,seq_loop_csv_dumper_235);
    seq_loop_csv_dumper_236 = new("./seq_loop_status236.csv");
    seq_loop_monitor_236 = new(seq_loop_intf_236,seq_loop_csv_dumper_236);
    seq_loop_csv_dumper_237 = new("./seq_loop_status237.csv");
    seq_loop_monitor_237 = new(seq_loop_intf_237,seq_loop_csv_dumper_237);
    seq_loop_csv_dumper_238 = new("./seq_loop_status238.csv");
    seq_loop_monitor_238 = new(seq_loop_intf_238,seq_loop_csv_dumper_238);
    seq_loop_csv_dumper_239 = new("./seq_loop_status239.csv");
    seq_loop_monitor_239 = new(seq_loop_intf_239,seq_loop_csv_dumper_239);
    seq_loop_csv_dumper_240 = new("./seq_loop_status240.csv");
    seq_loop_monitor_240 = new(seq_loop_intf_240,seq_loop_csv_dumper_240);
    seq_loop_csv_dumper_241 = new("./seq_loop_status241.csv");
    seq_loop_monitor_241 = new(seq_loop_intf_241,seq_loop_csv_dumper_241);
    seq_loop_csv_dumper_242 = new("./seq_loop_status242.csv");
    seq_loop_monitor_242 = new(seq_loop_intf_242,seq_loop_csv_dumper_242);
    seq_loop_csv_dumper_243 = new("./seq_loop_status243.csv");
    seq_loop_monitor_243 = new(seq_loop_intf_243,seq_loop_csv_dumper_243);
    seq_loop_csv_dumper_244 = new("./seq_loop_status244.csv");
    seq_loop_monitor_244 = new(seq_loop_intf_244,seq_loop_csv_dumper_244);
    seq_loop_csv_dumper_245 = new("./seq_loop_status245.csv");
    seq_loop_monitor_245 = new(seq_loop_intf_245,seq_loop_csv_dumper_245);
    seq_loop_csv_dumper_246 = new("./seq_loop_status246.csv");
    seq_loop_monitor_246 = new(seq_loop_intf_246,seq_loop_csv_dumper_246);
    seq_loop_csv_dumper_247 = new("./seq_loop_status247.csv");
    seq_loop_monitor_247 = new(seq_loop_intf_247,seq_loop_csv_dumper_247);
    seq_loop_csv_dumper_248 = new("./seq_loop_status248.csv");
    seq_loop_monitor_248 = new(seq_loop_intf_248,seq_loop_csv_dumper_248);
    seq_loop_csv_dumper_249 = new("./seq_loop_status249.csv");
    seq_loop_monitor_249 = new(seq_loop_intf_249,seq_loop_csv_dumper_249);
    seq_loop_csv_dumper_250 = new("./seq_loop_status250.csv");
    seq_loop_monitor_250 = new(seq_loop_intf_250,seq_loop_csv_dumper_250);
    seq_loop_csv_dumper_251 = new("./seq_loop_status251.csv");
    seq_loop_monitor_251 = new(seq_loop_intf_251,seq_loop_csv_dumper_251);
    seq_loop_csv_dumper_252 = new("./seq_loop_status252.csv");
    seq_loop_monitor_252 = new(seq_loop_intf_252,seq_loop_csv_dumper_252);
    seq_loop_csv_dumper_253 = new("./seq_loop_status253.csv");
    seq_loop_monitor_253 = new(seq_loop_intf_253,seq_loop_csv_dumper_253);


    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(module_monitor_7);
    sample_manager_inst.add_one_monitor(module_monitor_8);
    sample_manager_inst.add_one_monitor(module_monitor_9);
    sample_manager_inst.add_one_monitor(module_monitor_10);
    sample_manager_inst.add_one_monitor(module_monitor_11);
    sample_manager_inst.add_one_monitor(module_monitor_12);
    sample_manager_inst.add_one_monitor(module_monitor_13);
    sample_manager_inst.add_one_monitor(module_monitor_14);
    sample_manager_inst.add_one_monitor(module_monitor_15);
    sample_manager_inst.add_one_monitor(module_monitor_16);
    sample_manager_inst.add_one_monitor(module_monitor_17);
    sample_manager_inst.add_one_monitor(module_monitor_18);
    sample_manager_inst.add_one_monitor(module_monitor_19);
    sample_manager_inst.add_one_monitor(module_monitor_20);
    sample_manager_inst.add_one_monitor(module_monitor_21);
    sample_manager_inst.add_one_monitor(module_monitor_22);
    sample_manager_inst.add_one_monitor(module_monitor_23);
    sample_manager_inst.add_one_monitor(module_monitor_24);
    sample_manager_inst.add_one_monitor(module_monitor_25);
    sample_manager_inst.add_one_monitor(module_monitor_26);
    sample_manager_inst.add_one_monitor(module_monitor_27);
    sample_manager_inst.add_one_monitor(module_monitor_28);
    sample_manager_inst.add_one_monitor(module_monitor_29);
    sample_manager_inst.add_one_monitor(module_monitor_30);
    sample_manager_inst.add_one_monitor(module_monitor_31);
    sample_manager_inst.add_one_monitor(module_monitor_32);
    sample_manager_inst.add_one_monitor(module_monitor_33);
    sample_manager_inst.add_one_monitor(module_monitor_34);
    sample_manager_inst.add_one_monitor(module_monitor_35);
    sample_manager_inst.add_one_monitor(module_monitor_36);
    sample_manager_inst.add_one_monitor(module_monitor_37);
    sample_manager_inst.add_one_monitor(module_monitor_38);
    sample_manager_inst.add_one_monitor(module_monitor_39);
    sample_manager_inst.add_one_monitor(module_monitor_40);
    sample_manager_inst.add_one_monitor(module_monitor_41);
    sample_manager_inst.add_one_monitor(module_monitor_42);
    sample_manager_inst.add_one_monitor(module_monitor_43);
    sample_manager_inst.add_one_monitor(module_monitor_44);
    sample_manager_inst.add_one_monitor(module_monitor_45);
    sample_manager_inst.add_one_monitor(module_monitor_46);
    sample_manager_inst.add_one_monitor(module_monitor_47);
    sample_manager_inst.add_one_monitor(module_monitor_48);
    sample_manager_inst.add_one_monitor(module_monitor_49);
    sample_manager_inst.add_one_monitor(module_monitor_50);
    sample_manager_inst.add_one_monitor(module_monitor_51);
    sample_manager_inst.add_one_monitor(module_monitor_52);
    sample_manager_inst.add_one_monitor(module_monitor_53);
    sample_manager_inst.add_one_monitor(module_monitor_54);
    sample_manager_inst.add_one_monitor(module_monitor_55);
    sample_manager_inst.add_one_monitor(module_monitor_56);
    sample_manager_inst.add_one_monitor(module_monitor_57);
    sample_manager_inst.add_one_monitor(module_monitor_58);
    sample_manager_inst.add_one_monitor(module_monitor_59);
    sample_manager_inst.add_one_monitor(module_monitor_60);
    sample_manager_inst.add_one_monitor(module_monitor_61);
    sample_manager_inst.add_one_monitor(module_monitor_62);
    sample_manager_inst.add_one_monitor(module_monitor_63);
    sample_manager_inst.add_one_monitor(module_monitor_64);
    sample_manager_inst.add_one_monitor(module_monitor_65);
    sample_manager_inst.add_one_monitor(module_monitor_66);
    sample_manager_inst.add_one_monitor(module_monitor_67);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_7);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_8);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_9);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_10);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_11);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_12);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_13);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_14);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_15);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_16);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_17);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_18);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_19);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_20);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_21);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_22);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_23);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_24);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_25);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_26);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_27);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_28);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_29);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_30);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_31);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_32);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_33);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_34);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_35);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_36);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_37);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_38);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_39);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_40);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_41);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_42);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_43);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_44);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_45);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_46);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_47);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_48);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_49);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_50);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_51);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_52);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_53);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_54);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_55);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_56);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_57);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_58);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_59);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_60);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_61);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_62);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_63);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_64);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_65);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_66);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_67);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_68);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_69);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_70);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_71);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_72);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_73);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_74);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_75);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_76);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_77);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_78);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_79);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_80);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_81);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_82);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_83);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_84);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_85);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_86);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_87);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_88);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_89);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_90);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_91);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_92);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_93);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_94);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_95);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_96);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_97);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_98);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_99);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_100);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_101);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_102);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_103);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_104);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_105);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_106);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_107);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_108);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_109);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_110);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_111);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_112);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_113);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_114);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_115);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_116);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_117);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_118);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_119);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_120);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_121);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_122);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_123);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_124);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_125);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_126);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_127);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_128);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_129);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_130);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_131);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_132);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_133);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_134);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_135);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_136);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_137);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_138);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_139);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_140);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_141);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_142);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_143);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_144);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_145);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_146);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_147);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_148);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_149);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_150);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_151);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_152);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_153);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_154);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_155);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_156);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_157);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_158);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_159);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_160);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_161);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_162);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_163);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_164);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_165);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_166);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_167);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_168);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_169);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_170);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_171);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_172);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_173);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_174);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_175);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_176);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_177);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_178);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_179);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_180);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_181);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_182);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_183);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_184);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_185);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_186);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_187);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_188);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_189);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_190);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_191);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_192);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_193);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_194);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_195);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_196);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_197);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_198);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_199);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_200);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_201);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_202);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_203);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_204);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_205);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_206);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_207);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_208);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_209);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_210);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_211);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_212);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_213);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_214);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_215);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_216);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_217);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_218);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_219);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_220);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_221);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_222);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_223);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_224);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_225);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_226);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_227);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_228);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_229);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_230);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_231);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_232);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_233);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_234);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_235);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_236);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_237);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_238);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_239);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_240);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_241);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_242);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_243);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_244);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_245);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_246);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_247);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_248);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_249);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_250);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_251);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_252);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_253);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1) begin
                @(negedge clock);
                break;
            end
            else
                @(posedge clock);
        end
    endtask


endmodule
